
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_router_pl is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type UNSIGNED is array (INTEGER range <>) of std_logic;
subtype vc_status_vec is std_logic_vector (1 downto 0);
type vc_status_array is array (INTEGER range <>) of vc_status_vec;
subtype vc_status_vec_enc is std_logic_vector (0 downto 0);
type vc_status_array_enc is array (INTEGER range <>) of vc_status_vec_enc;
subtype flit is std_logic_vector (63 downto 0);
type VHDLOUT_TYPE is array (0 downto 0) of std_logic_vector (9 downto 0);
type VHDLOUT_TYPE_2 is array (12 downto 0) of std_logic_vector (9 downto 0);
type flit_vector is array (INTEGER range <>) of std_logic_vector (63 downto 0);

end CONV_PACK_router_pl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity switch_allocator_7_DXYU_DW_mod_tc_6 is

   port( a : in std_logic_vector (4 downto 0);  b : in std_logic_vector (31 
         downto 0);  quotient : out std_logic_vector (4 downto 0);  remainder :
         out std_logic_vector (31 downto 0);  divide_by_0 : out std_logic);

end switch_allocator_7_DXYU_DW_mod_tc_6;

architecture SYN_cla of switch_allocator_7_DXYU_DW_mod_tc_6 is

   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22xp33_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp33_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND5xp2_ASAP7_75t_R
      port( A, B, C, D, E : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal u_div_MAdd_0_port, u_div_MAdd_1_port, u_div_MAdd_2_port, 
      u_div_SumTmp_0_1_port, u_div_SumTmp_0_2_port, u_div_SumTmp_0_3_port, 
      u_div_SumTmp_0_4_port, u_div_SumTmp_1_1_port, u_div_SumTmp_1_2_port, 
      u_div_CryTmp_0_5_port, u_div_CryTmp_1_4_port, u_div_PartRem_1_1_port, 
      u_div_PartRem_1_2_port, u_div_PartRem_1_3_port, u_div_PartRem_1_4_port, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18 : std_logic;

begin
   
   U1 : NOR2xp33_ASAP7_75t_R port map( A => n11, B => n6, Y => 
                           u_div_CryTmp_1_4_port);
   U2 : NOR2xp33_ASAP7_75t_R port map( A => n5, B => n12, Y => 
                           u_div_PartRem_1_4_port);
   U3 : INVx1_ASAP7_75t_R port map( A => a(0), Y => n1);
   U4 : INVx1_ASAP7_75t_R port map( A => n16, Y => u_div_MAdd_1_port);
   U5 : INVx1_ASAP7_75t_R port map( A => n17, Y => u_div_MAdd_0_port);
   U6 : INVx1_ASAP7_75t_R port map( A => n15, Y => u_div_MAdd_2_port);
   U7 : INVx1_ASAP7_75t_R port map( A => u_div_CryTmp_0_5_port, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => u_div_PartRem_1_2_port, Y => n3);
   U9 : INVx1_ASAP7_75t_R port map( A => u_div_PartRem_1_3_port, Y => n4);
   U10 : INVx1_ASAP7_75t_R port map( A => u_div_CryTmp_1_4_port, Y => n5);
   U11 : INVx1_ASAP7_75t_R port map( A => a(3), Y => n6);
   U12 : INVx1_ASAP7_75t_R port map( A => a(1), Y => n7);
   U13 : NAND2xp33_ASAP7_75t_R port map( A => a(0), B => u_div_PartRem_1_1_port
                           , Y => n8);
   U14 : AOI22xp33_ASAP7_75t_R port map( A1 => n8, A2 => n4, B1 => n3, B2 => n4
                           , Y => n10);
   U15 : OR2x2_ASAP7_75t_R port map( A => n10, B => u_div_PartRem_1_4_port, Y 
                           => u_div_CryTmp_0_5_port);
   U16 : XOR2xp5_ASAP7_75t_R port map( A => a(0), B => u_div_PartRem_1_1_port, 
                           Y => u_div_SumTmp_0_1_port);
   U17 : XNOR2xp5_ASAP7_75t_R port map( A => u_div_PartRem_1_2_port, B => n8, Y
                           => u_div_SumTmp_0_2_port);
   U18 : NOR2xp33_ASAP7_75t_R port map( A => n8, B => n3, Y => n9);
   U19 : XNOR2xp5_ASAP7_75t_R port map( A => u_div_PartRem_1_3_port, B => n9, Y
                           => u_div_SumTmp_0_3_port);
   U20 : XNOR2xp5_ASAP7_75t_R port map( A => u_div_PartRem_1_4_port, B => n10, 
                           Y => u_div_SumTmp_0_4_port);
   U21 : NAND2xp33_ASAP7_75t_R port map( A => a(1), B => a(2), Y => n11);
   U22 : XOR2xp5_ASAP7_75t_R port map( A => a(1), B => a(2), Y => 
                           u_div_SumTmp_1_1_port);
   U23 : XOR2xp5_ASAP7_75t_R port map( A => n6, B => n11, Y => 
                           u_div_SumTmp_1_2_port);
   U24 : NOR2xp33_ASAP7_75t_R port map( A => n11, B => n6, Y => n12);
   U25 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_2_port, B => n18, Y => 
                           remainder(2));
   U26 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_1_port, B => n18, Y => 
                           remainder(1));
   U27 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_0_port, B => n18, Y => 
                           remainder(0));
   U28 : NAND5xp2_ASAP7_75t_R port map( A => n14, B => n13, C => n15, D => n17,
                           E => n16, Y => n18);
   U29 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_1_port, A2 => 
                           u_div_CryTmp_0_5_port, B1 => u_div_PartRem_1_1_port,
                           B2 => n2, Y => n16);
   U30 : OAI22xp33_ASAP7_75t_R port map( A1 => a(1), A2 => n5, B1 => 
                           u_div_CryTmp_1_4_port, B2 => n7, Y => 
                           u_div_PartRem_1_1_port);
   U31 : AOI22xp33_ASAP7_75t_R port map( A1 => n1, A2 => u_div_CryTmp_0_5_port,
                           B1 => n2, B2 => a(0), Y => n17);
   U32 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_2_port, A2 => 
                           u_div_CryTmp_0_5_port, B1 => u_div_PartRem_1_2_port,
                           B2 => n2, Y => n15);
   U33 : AO22x1_ASAP7_75t_R port map( A1 => u_div_SumTmp_1_1_port, A2 => 
                           u_div_CryTmp_1_4_port, B1 => a(2), B2 => n5, Y => 
                           u_div_PartRem_1_2_port);
   U34 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_4_port, A2 => 
                           u_div_CryTmp_0_5_port, B1 => u_div_PartRem_1_4_port,
                           B2 => n2, Y => n13);
   U35 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_3_port, A2 => 
                           u_div_CryTmp_0_5_port, B1 => u_div_PartRem_1_3_port,
                           B2 => n2, Y => n14);
   U36 : AO22x1_ASAP7_75t_R port map( A1 => u_div_SumTmp_1_2_port, A2 => 
                           u_div_CryTmp_1_4_port, B1 => a(3), B2 => n5, Y => 
                           u_div_PartRem_1_3_port);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity switch_allocator_7_DXYU_DW_mod_tc_5 is

   port( a : in std_logic_vector (5 downto 0);  b : in std_logic_vector (31 
         downto 0);  quotient : out std_logic_vector (5 downto 0);  remainder :
         out std_logic_vector (31 downto 0);  divide_by_0 : out std_logic);

end switch_allocator_7_DXYU_DW_mod_tc_5;

architecture SYN_cla of switch_allocator_7_DXYU_DW_mod_tc_5 is

   component AOI22xp33_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp33_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AND3x1_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal u_div_MAdd_0_port, u_div_MAdd_1_port, u_div_MAdd_2_port, 
      u_div_SumTmp_0_1_port, u_div_SumTmp_0_2_port, u_div_SumTmp_0_3_port, 
      u_div_SumTmp_0_4_port, u_div_SumTmp_1_1_port, u_div_SumTmp_1_2_port, 
      u_div_CryTmp_0_6_port, u_div_CryTmp_1_5_port, u_div_PartRem_1_1_port, 
      u_div_PartRem_1_2_port, u_div_PartRem_1_3_port, u_div_PartRem_1_4_port, 
      u_div_u_add_PartRem_3_0_SUM_4_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n6, Y => 
                           u_div_CryTmp_1_5_port);
   U2 : NOR2xp33_ASAP7_75t_R port map( A => n5, B => n10, Y => 
                           u_div_PartRem_1_4_port);
   U3 : NAND2xp33_ASAP7_75t_R port map( A => a(0), B => u_div_PartRem_1_1_port,
                           Y => n1);
   U4 : NOR2xp33_ASAP7_75t_R port map( A => n4, B => n1, Y => n2);
   U5 : OR2x2_ASAP7_75t_R port map( A => u_div_PartRem_1_3_port, B => n2, Y => 
                           n3);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => n3, B => u_div_PartRem_1_4_port, Y 
                           => u_div_u_add_PartRem_3_0_SUM_4_port);
   U7 : XOR2xp5_ASAP7_75t_R port map( A => a(0), B => u_div_PartRem_1_1_port, Y
                           => u_div_SumTmp_0_1_port);
   U8 : XOR2xp5_ASAP7_75t_R port map( A => n4, B => n1, Y => 
                           u_div_SumTmp_0_2_port);
   U9 : XNOR2xp5_ASAP7_75t_R port map( A => u_div_PartRem_1_3_port, B => n2, Y 
                           => u_div_SumTmp_0_3_port);
   U10 : XNOR2xp5_ASAP7_75t_R port map( A => u_div_PartRem_1_4_port, B => n3, Y
                           => u_div_SumTmp_0_4_port);
   U11 : INVx1_ASAP7_75t_R port map( A => u_div_PartRem_1_2_port, Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => u_div_u_add_PartRem_3_0_SUM_4_port, Y
                           => u_div_CryTmp_0_6_port);
   U13 : INVx1_ASAP7_75t_R port map( A => n14, Y => u_div_MAdd_1_port);
   U14 : INVx1_ASAP7_75t_R port map( A => n13, Y => u_div_MAdd_2_port);
   U15 : INVx1_ASAP7_75t_R port map( A => n15, Y => u_div_MAdd_0_port);
   U16 : INVx1_ASAP7_75t_R port map( A => u_div_CryTmp_1_5_port, Y => n5);
   U17 : INVx1_ASAP7_75t_R port map( A => a(3), Y => n6);
   U18 : INVx1_ASAP7_75t_R port map( A => a(1), Y => n7);
   U19 : INVx1_ASAP7_75t_R port map( A => a(0), Y => n8);
   U20 : NAND3xp33_ASAP7_75t_R port map( A => n12, B => n17, C => n11, Y => n16
                           );
   U21 : NAND2xp33_ASAP7_75t_R port map( A => a(1), B => a(2), Y => n9);
   U22 : XOR2xp5_ASAP7_75t_R port map( A => a(1), B => a(2), Y => 
                           u_div_SumTmp_1_1_port);
   U23 : XNOR2xp5_ASAP7_75t_R port map( A => a(3), B => n9, Y => 
                           u_div_SumTmp_1_2_port);
   U24 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n6, Y => n10);
   U25 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_2_port, B => n16, Y => 
                           remainder(2));
   U26 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_1_port, B => n16, Y => 
                           remainder(1));
   U27 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_0_port, B => n16, Y => 
                           remainder(0));
   U28 : AND3x1_ASAP7_75t_R port map( A => n15, B => n13, C => n14, Y => n17);
   U29 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_1_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_1_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n14);
   U30 : OAI22xp33_ASAP7_75t_R port map( A1 => a(1), A2 => n5, B1 => 
                           u_div_CryTmp_1_5_port, B2 => n7, Y => 
                           u_div_PartRem_1_1_port);
   U31 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_2_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_2_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n13);
   U32 : AO22x1_ASAP7_75t_R port map( A1 => u_div_SumTmp_1_1_port, A2 => 
                           u_div_CryTmp_1_5_port, B1 => a(2), B2 => n5, Y => 
                           u_div_PartRem_1_2_port);
   U33 : AOI22xp33_ASAP7_75t_R port map( A1 => n8, A2 => u_div_CryTmp_0_6_port,
                           B1 => u_div_u_add_PartRem_3_0_SUM_4_port, B2 => a(0)
                           , Y => n15);
   U34 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_3_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_3_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n12);
   U35 : AO22x1_ASAP7_75t_R port map( A1 => u_div_SumTmp_1_2_port, A2 => 
                           u_div_CryTmp_1_5_port, B1 => a(3), B2 => n5, Y => 
                           u_div_PartRem_1_3_port);
   U36 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_4_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_4_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n11);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity switch_allocator_7_DXYU_DW_mod_tc_4 is

   port( a : in std_logic_vector (5 downto 0);  b : in std_logic_vector (31 
         downto 0);  quotient : out std_logic_vector (5 downto 0);  remainder :
         out std_logic_vector (31 downto 0);  divide_by_0 : out std_logic);

end switch_allocator_7_DXYU_DW_mod_tc_4;

architecture SYN_cla of switch_allocator_7_DXYU_DW_mod_tc_4 is

   component AOI22xp33_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp33_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AND3x1_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal u_div_MAdd_0_port, u_div_MAdd_1_port, u_div_MAdd_2_port, 
      u_div_SumTmp_0_1_port, u_div_SumTmp_0_2_port, u_div_SumTmp_0_3_port, 
      u_div_SumTmp_0_4_port, u_div_SumTmp_1_1_port, u_div_SumTmp_1_2_port, 
      u_div_CryTmp_0_6_port, u_div_CryTmp_1_5_port, u_div_PartRem_1_1_port, 
      u_div_PartRem_1_2_port, u_div_PartRem_1_3_port, u_div_PartRem_1_4_port, 
      u_div_u_add_PartRem_3_0_SUM_4_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n6, Y => 
                           u_div_CryTmp_1_5_port);
   U2 : NOR2xp33_ASAP7_75t_R port map( A => n5, B => n10, Y => 
                           u_div_PartRem_1_4_port);
   U3 : NAND2xp33_ASAP7_75t_R port map( A => a(0), B => u_div_PartRem_1_1_port,
                           Y => n1);
   U4 : NOR2xp33_ASAP7_75t_R port map( A => n4, B => n1, Y => n2);
   U5 : OR2x2_ASAP7_75t_R port map( A => u_div_PartRem_1_3_port, B => n2, Y => 
                           n3);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => n3, B => u_div_PartRem_1_4_port, Y 
                           => u_div_u_add_PartRem_3_0_SUM_4_port);
   U7 : XOR2xp5_ASAP7_75t_R port map( A => a(0), B => u_div_PartRem_1_1_port, Y
                           => u_div_SumTmp_0_1_port);
   U8 : XOR2xp5_ASAP7_75t_R port map( A => n4, B => n1, Y => 
                           u_div_SumTmp_0_2_port);
   U9 : XNOR2xp5_ASAP7_75t_R port map( A => u_div_PartRem_1_3_port, B => n2, Y 
                           => u_div_SumTmp_0_3_port);
   U10 : XNOR2xp5_ASAP7_75t_R port map( A => u_div_PartRem_1_4_port, B => n3, Y
                           => u_div_SumTmp_0_4_port);
   U11 : INVx1_ASAP7_75t_R port map( A => u_div_PartRem_1_2_port, Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => u_div_u_add_PartRem_3_0_SUM_4_port, Y
                           => u_div_CryTmp_0_6_port);
   U13 : INVx1_ASAP7_75t_R port map( A => n14, Y => u_div_MAdd_1_port);
   U14 : INVx1_ASAP7_75t_R port map( A => n13, Y => u_div_MAdd_2_port);
   U15 : INVx1_ASAP7_75t_R port map( A => n15, Y => u_div_MAdd_0_port);
   U16 : INVx1_ASAP7_75t_R port map( A => u_div_CryTmp_1_5_port, Y => n5);
   U17 : INVx1_ASAP7_75t_R port map( A => a(3), Y => n6);
   U18 : INVx1_ASAP7_75t_R port map( A => a(1), Y => n7);
   U19 : INVx1_ASAP7_75t_R port map( A => a(0), Y => n8);
   U20 : NAND3xp33_ASAP7_75t_R port map( A => n12, B => n17, C => n11, Y => n16
                           );
   U21 : NAND2xp33_ASAP7_75t_R port map( A => a(1), B => a(2), Y => n9);
   U22 : XOR2xp5_ASAP7_75t_R port map( A => a(1), B => a(2), Y => 
                           u_div_SumTmp_1_1_port);
   U23 : XNOR2xp5_ASAP7_75t_R port map( A => a(3), B => n9, Y => 
                           u_div_SumTmp_1_2_port);
   U24 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n6, Y => n10);
   U25 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_2_port, B => n16, Y => 
                           remainder(2));
   U26 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_1_port, B => n16, Y => 
                           remainder(1));
   U27 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_0_port, B => n16, Y => 
                           remainder(0));
   U28 : AND3x1_ASAP7_75t_R port map( A => n15, B => n13, C => n14, Y => n17);
   U29 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_1_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_1_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n14);
   U30 : OAI22xp33_ASAP7_75t_R port map( A1 => a(1), A2 => n5, B1 => 
                           u_div_CryTmp_1_5_port, B2 => n7, Y => 
                           u_div_PartRem_1_1_port);
   U31 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_2_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_2_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n13);
   U32 : AO22x1_ASAP7_75t_R port map( A1 => u_div_SumTmp_1_1_port, A2 => 
                           u_div_CryTmp_1_5_port, B1 => a(2), B2 => n5, Y => 
                           u_div_PartRem_1_2_port);
   U33 : AOI22xp33_ASAP7_75t_R port map( A1 => n8, A2 => u_div_CryTmp_0_6_port,
                           B1 => u_div_u_add_PartRem_3_0_SUM_4_port, B2 => a(0)
                           , Y => n15);
   U34 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_3_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_3_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n12);
   U35 : AO22x1_ASAP7_75t_R port map( A1 => u_div_SumTmp_1_2_port, A2 => 
                           u_div_CryTmp_1_5_port, B1 => a(3), B2 => n5, Y => 
                           u_div_PartRem_1_3_port);
   U36 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_4_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_4_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n11);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity switch_allocator_7_DXYU_DW_mod_tc_3 is

   port( a : in std_logic_vector (5 downto 0);  b : in std_logic_vector (31 
         downto 0);  quotient : out std_logic_vector (5 downto 0);  remainder :
         out std_logic_vector (31 downto 0);  divide_by_0 : out std_logic);

end switch_allocator_7_DXYU_DW_mod_tc_3;

architecture SYN_cla of switch_allocator_7_DXYU_DW_mod_tc_3 is

   component AOI22xp33_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp33_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AND3x1_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal u_div_MAdd_0_port, u_div_MAdd_1_port, u_div_MAdd_2_port, 
      u_div_SumTmp_0_1_port, u_div_SumTmp_0_2_port, u_div_SumTmp_0_3_port, 
      u_div_SumTmp_0_4_port, u_div_SumTmp_1_1_port, u_div_SumTmp_1_2_port, 
      u_div_CryTmp_0_6_port, u_div_CryTmp_1_5_port, u_div_PartRem_1_1_port, 
      u_div_PartRem_1_2_port, u_div_PartRem_1_3_port, u_div_PartRem_1_4_port, 
      u_div_u_add_PartRem_3_0_SUM_4_port, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => a(2), Y => 
                           u_div_CryTmp_1_5_port);
   U2 : NOR2xp33_ASAP7_75t_R port map( A => n6, B => n10, Y => 
                           u_div_PartRem_1_4_port);
   U3 : NAND2xp33_ASAP7_75t_R port map( A => a(0), B => u_div_PartRem_1_1_port,
                           Y => n2);
   U4 : NOR2xp33_ASAP7_75t_R port map( A => n5, B => n2, Y => n3);
   U5 : OR2x2_ASAP7_75t_R port map( A => u_div_PartRem_1_3_port, B => n3, Y => 
                           n4);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => n4, B => u_div_PartRem_1_4_port, Y 
                           => u_div_u_add_PartRem_3_0_SUM_4_port);
   U7 : XOR2xp5_ASAP7_75t_R port map( A => a(0), B => u_div_PartRem_1_1_port, Y
                           => u_div_SumTmp_0_1_port);
   U8 : XOR2xp5_ASAP7_75t_R port map( A => n5, B => n2, Y => 
                           u_div_SumTmp_0_2_port);
   U9 : XNOR2xp5_ASAP7_75t_R port map( A => u_div_PartRem_1_3_port, B => n3, Y 
                           => u_div_SumTmp_0_3_port);
   U10 : XNOR2xp5_ASAP7_75t_R port map( A => u_div_PartRem_1_4_port, B => n4, Y
                           => u_div_SumTmp_0_4_port);
   U11 : INVx1_ASAP7_75t_R port map( A => u_div_PartRem_1_2_port, Y => n5);
   U12 : INVx1_ASAP7_75t_R port map( A => u_div_u_add_PartRem_3_0_SUM_4_port, Y
                           => u_div_CryTmp_0_6_port);
   U13 : INVx1_ASAP7_75t_R port map( A => n14, Y => u_div_MAdd_1_port);
   U14 : INVx1_ASAP7_75t_R port map( A => n13, Y => u_div_MAdd_2_port);
   U15 : INVx1_ASAP7_75t_R port map( A => n15, Y => u_div_MAdd_0_port);
   U16 : INVx1_ASAP7_75t_R port map( A => u_div_CryTmp_1_5_port, Y => n6);
   U17 : INVx1_ASAP7_75t_R port map( A => a(1), Y => n7);
   U18 : INVx1_ASAP7_75t_R port map( A => a(0), Y => n8);
   U19 : NAND3xp33_ASAP7_75t_R port map( A => n12, B => n17, C => n11, Y => n16
                           );
   U20 : NAND2xp33_ASAP7_75t_R port map( A => a(1), B => a(2), Y => n9);
   U21 : XOR2xp5_ASAP7_75t_R port map( A => a(1), B => a(2), Y => 
                           u_div_SumTmp_1_1_port);
   U22 : XNOR2xp5_ASAP7_75t_R port map( A => a(3), B => n9, Y => 
                           u_div_SumTmp_1_2_port);
   U23 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => a(2), Y => n10);
   U24 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_2_port, B => n16, Y => 
                           remainder(2));
   U25 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_1_port, B => n16, Y => 
                           remainder(1));
   U26 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_0_port, B => n16, Y => 
                           remainder(0));
   U27 : AND3x1_ASAP7_75t_R port map( A => n15, B => n13, C => n14, Y => n17);
   U28 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_1_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_1_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n14);
   U29 : OAI22xp33_ASAP7_75t_R port map( A1 => a(1), A2 => n6, B1 => 
                           u_div_CryTmp_1_5_port, B2 => n7, Y => 
                           u_div_PartRem_1_1_port);
   U30 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_2_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_2_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n13);
   U31 : AO22x1_ASAP7_75t_R port map( A1 => u_div_SumTmp_1_1_port, A2 => 
                           u_div_CryTmp_1_5_port, B1 => a(2), B2 => n6, Y => 
                           u_div_PartRem_1_2_port);
   U32 : AOI22xp33_ASAP7_75t_R port map( A1 => n8, A2 => u_div_CryTmp_0_6_port,
                           B1 => u_div_u_add_PartRem_3_0_SUM_4_port, B2 => a(0)
                           , Y => n15);
   U33 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_3_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_3_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n12);
   U34 : AO22x1_ASAP7_75t_R port map( A1 => u_div_SumTmp_1_2_port, A2 => 
                           u_div_CryTmp_1_5_port, B1 => a(3), B2 => n6, Y => 
                           u_div_PartRem_1_3_port);
   U35 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_4_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_4_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n11);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity switch_allocator_7_DXYU_DW_mod_tc_2 is

   port( a : in std_logic_vector (5 downto 0);  b : in std_logic_vector (31 
         downto 0);  quotient : out std_logic_vector (5 downto 0);  remainder :
         out std_logic_vector (31 downto 0);  divide_by_0 : out std_logic);

end switch_allocator_7_DXYU_DW_mod_tc_2;

architecture SYN_cla of switch_allocator_7_DXYU_DW_mod_tc_2 is

   component AOI22xp33_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp33_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AND3x1_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal u_div_MAdd_0_port, u_div_MAdd_1_port, u_div_MAdd_2_port, 
      u_div_SumTmp_0_1_port, u_div_SumTmp_0_2_port, u_div_SumTmp_0_3_port, 
      u_div_SumTmp_0_4_port, u_div_SumTmp_1_1_port, u_div_SumTmp_1_2_port, 
      u_div_CryTmp_0_6_port, u_div_CryTmp_1_5_port, u_div_PartRem_1_1_port, 
      u_div_PartRem_1_2_port, u_div_PartRem_1_3_port, u_div_PartRem_1_4_port, 
      u_div_u_add_PartRem_3_0_SUM_4_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n6, Y => 
                           u_div_CryTmp_1_5_port);
   U2 : NOR2xp33_ASAP7_75t_R port map( A => n5, B => n10, Y => 
                           u_div_PartRem_1_4_port);
   U3 : NAND2xp33_ASAP7_75t_R port map( A => a(0), B => u_div_PartRem_1_1_port,
                           Y => n1);
   U4 : NOR2xp33_ASAP7_75t_R port map( A => n4, B => n1, Y => n2);
   U5 : OR2x2_ASAP7_75t_R port map( A => u_div_PartRem_1_3_port, B => n2, Y => 
                           n3);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => n3, B => u_div_PartRem_1_4_port, Y 
                           => u_div_u_add_PartRem_3_0_SUM_4_port);
   U7 : XOR2xp5_ASAP7_75t_R port map( A => a(0), B => u_div_PartRem_1_1_port, Y
                           => u_div_SumTmp_0_1_port);
   U8 : XOR2xp5_ASAP7_75t_R port map( A => n4, B => n1, Y => 
                           u_div_SumTmp_0_2_port);
   U9 : XNOR2xp5_ASAP7_75t_R port map( A => u_div_PartRem_1_3_port, B => n2, Y 
                           => u_div_SumTmp_0_3_port);
   U10 : XNOR2xp5_ASAP7_75t_R port map( A => u_div_PartRem_1_4_port, B => n3, Y
                           => u_div_SumTmp_0_4_port);
   U11 : INVx1_ASAP7_75t_R port map( A => u_div_PartRem_1_2_port, Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => u_div_u_add_PartRem_3_0_SUM_4_port, Y
                           => u_div_CryTmp_0_6_port);
   U13 : INVx1_ASAP7_75t_R port map( A => n14, Y => u_div_MAdd_1_port);
   U14 : INVx1_ASAP7_75t_R port map( A => n13, Y => u_div_MAdd_2_port);
   U15 : INVx1_ASAP7_75t_R port map( A => n15, Y => u_div_MAdd_0_port);
   U16 : INVx1_ASAP7_75t_R port map( A => u_div_CryTmp_1_5_port, Y => n5);
   U17 : INVx1_ASAP7_75t_R port map( A => a(3), Y => n6);
   U18 : INVx1_ASAP7_75t_R port map( A => a(1), Y => n7);
   U19 : INVx1_ASAP7_75t_R port map( A => a(0), Y => n8);
   U20 : NAND3xp33_ASAP7_75t_R port map( A => n12, B => n17, C => n11, Y => n16
                           );
   U21 : NAND2xp33_ASAP7_75t_R port map( A => a(1), B => a(2), Y => n9);
   U22 : XOR2xp5_ASAP7_75t_R port map( A => a(1), B => a(2), Y => 
                           u_div_SumTmp_1_1_port);
   U23 : XNOR2xp5_ASAP7_75t_R port map( A => a(3), B => n9, Y => 
                           u_div_SumTmp_1_2_port);
   U24 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n6, Y => n10);
   U25 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_2_port, B => n16, Y => 
                           remainder(2));
   U26 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_1_port, B => n16, Y => 
                           remainder(1));
   U27 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_0_port, B => n16, Y => 
                           remainder(0));
   U28 : AND3x1_ASAP7_75t_R port map( A => n15, B => n13, C => n14, Y => n17);
   U29 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_1_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_1_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n14);
   U30 : OAI22xp33_ASAP7_75t_R port map( A1 => a(1), A2 => n5, B1 => 
                           u_div_CryTmp_1_5_port, B2 => n7, Y => 
                           u_div_PartRem_1_1_port);
   U31 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_2_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_2_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n13);
   U32 : AO22x1_ASAP7_75t_R port map( A1 => u_div_SumTmp_1_1_port, A2 => 
                           u_div_CryTmp_1_5_port, B1 => a(2), B2 => n5, Y => 
                           u_div_PartRem_1_2_port);
   U33 : AOI22xp33_ASAP7_75t_R port map( A1 => n8, A2 => u_div_CryTmp_0_6_port,
                           B1 => u_div_u_add_PartRem_3_0_SUM_4_port, B2 => a(0)
                           , Y => n15);
   U34 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_3_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_3_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n12);
   U35 : AO22x1_ASAP7_75t_R port map( A1 => u_div_SumTmp_1_2_port, A2 => 
                           u_div_CryTmp_1_5_port, B1 => a(3), B2 => n5, Y => 
                           u_div_PartRem_1_3_port);
   U36 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_4_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_4_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n11);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity switch_allocator_7_DXYU_DW_mod_tc_1 is

   port( a : in std_logic_vector (5 downto 0);  b : in std_logic_vector (31 
         downto 0);  quotient : out std_logic_vector (5 downto 0);  remainder :
         out std_logic_vector (31 downto 0);  divide_by_0 : out std_logic);

end switch_allocator_7_DXYU_DW_mod_tc_1;

architecture SYN_cla of switch_allocator_7_DXYU_DW_mod_tc_1 is

   component AOI22xp33_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp33_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AND3x1_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal u_div_MAdd_0_port, u_div_MAdd_1_port, u_div_MAdd_2_port, 
      u_div_SumTmp_0_1_port, u_div_SumTmp_0_2_port, u_div_SumTmp_0_3_port, 
      u_div_SumTmp_0_4_port, u_div_SumTmp_1_1_port, u_div_SumTmp_1_2_port, 
      u_div_CryTmp_0_6_port, u_div_CryTmp_1_5_port, u_div_PartRem_1_1_port, 
      u_div_PartRem_1_2_port, u_div_PartRem_1_3_port, u_div_PartRem_1_4_port, 
      u_div_u_add_PartRem_3_0_SUM_4_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n6, Y => 
                           u_div_CryTmp_1_5_port);
   U2 : NOR2xp33_ASAP7_75t_R port map( A => n5, B => n10, Y => 
                           u_div_PartRem_1_4_port);
   U3 : NAND2xp33_ASAP7_75t_R port map( A => a(0), B => u_div_PartRem_1_1_port,
                           Y => n1);
   U4 : NOR2xp33_ASAP7_75t_R port map( A => n4, B => n1, Y => n2);
   U5 : OR2x2_ASAP7_75t_R port map( A => u_div_PartRem_1_3_port, B => n2, Y => 
                           n3);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => n3, B => u_div_PartRem_1_4_port, Y 
                           => u_div_u_add_PartRem_3_0_SUM_4_port);
   U7 : XOR2xp5_ASAP7_75t_R port map( A => a(0), B => u_div_PartRem_1_1_port, Y
                           => u_div_SumTmp_0_1_port);
   U8 : XOR2xp5_ASAP7_75t_R port map( A => n4, B => n1, Y => 
                           u_div_SumTmp_0_2_port);
   U9 : XNOR2xp5_ASAP7_75t_R port map( A => u_div_PartRem_1_3_port, B => n2, Y 
                           => u_div_SumTmp_0_3_port);
   U10 : XNOR2xp5_ASAP7_75t_R port map( A => u_div_PartRem_1_4_port, B => n3, Y
                           => u_div_SumTmp_0_4_port);
   U11 : INVx1_ASAP7_75t_R port map( A => u_div_PartRem_1_2_port, Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => u_div_u_add_PartRem_3_0_SUM_4_port, Y
                           => u_div_CryTmp_0_6_port);
   U13 : INVx1_ASAP7_75t_R port map( A => n14, Y => u_div_MAdd_1_port);
   U14 : INVx1_ASAP7_75t_R port map( A => n13, Y => u_div_MAdd_2_port);
   U15 : INVx1_ASAP7_75t_R port map( A => n15, Y => u_div_MAdd_0_port);
   U16 : INVx1_ASAP7_75t_R port map( A => u_div_CryTmp_1_5_port, Y => n5);
   U17 : INVx1_ASAP7_75t_R port map( A => a(3), Y => n6);
   U18 : INVx1_ASAP7_75t_R port map( A => a(1), Y => n7);
   U19 : INVx1_ASAP7_75t_R port map( A => a(0), Y => n8);
   U20 : NAND3xp33_ASAP7_75t_R port map( A => n12, B => n17, C => n11, Y => n16
                           );
   U21 : NAND2xp33_ASAP7_75t_R port map( A => a(1), B => a(2), Y => n9);
   U22 : XOR2xp5_ASAP7_75t_R port map( A => a(1), B => a(2), Y => 
                           u_div_SumTmp_1_1_port);
   U23 : XNOR2xp5_ASAP7_75t_R port map( A => a(3), B => n9, Y => 
                           u_div_SumTmp_1_2_port);
   U24 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n6, Y => n10);
   U25 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_2_port, B => n16, Y => 
                           remainder(2));
   U26 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_1_port, B => n16, Y => 
                           remainder(1));
   U27 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_0_port, B => n16, Y => 
                           remainder(0));
   U28 : AND3x1_ASAP7_75t_R port map( A => n15, B => n13, C => n14, Y => n17);
   U29 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_1_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_1_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n14);
   U30 : OAI22xp33_ASAP7_75t_R port map( A1 => a(1), A2 => n5, B1 => 
                           u_div_CryTmp_1_5_port, B2 => n7, Y => 
                           u_div_PartRem_1_1_port);
   U31 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_2_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_2_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n13);
   U32 : AO22x1_ASAP7_75t_R port map( A1 => u_div_SumTmp_1_1_port, A2 => 
                           u_div_CryTmp_1_5_port, B1 => a(2), B2 => n5, Y => 
                           u_div_PartRem_1_2_port);
   U33 : AOI22xp33_ASAP7_75t_R port map( A1 => n8, A2 => u_div_CryTmp_0_6_port,
                           B1 => u_div_u_add_PartRem_3_0_SUM_4_port, B2 => a(0)
                           , Y => n15);
   U34 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_3_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_3_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n12);
   U35 : AO22x1_ASAP7_75t_R port map( A1 => u_div_SumTmp_1_2_port, A2 => 
                           u_div_CryTmp_1_5_port, B1 => a(3), B2 => n5, Y => 
                           u_div_PartRem_1_3_port);
   U36 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_4_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_4_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n11);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity switch_allocator_7_DXYU_DW_mod_tc_0 is

   port( a : in std_logic_vector (5 downto 0);  b : in std_logic_vector (31 
         downto 0);  quotient : out std_logic_vector (5 downto 0);  remainder :
         out std_logic_vector (31 downto 0);  divide_by_0 : out std_logic);

end switch_allocator_7_DXYU_DW_mod_tc_0;

architecture SYN_cla of switch_allocator_7_DXYU_DW_mod_tc_0 is

   component AOI22xp33_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp33_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AND3x1_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal u_div_MAdd_0_port, u_div_MAdd_1_port, u_div_MAdd_2_port, 
      u_div_SumTmp_0_1_port, u_div_SumTmp_0_2_port, u_div_SumTmp_0_3_port, 
      u_div_SumTmp_0_4_port, u_div_SumTmp_1_1_port, u_div_SumTmp_1_2_port, 
      u_div_CryTmp_0_6_port, u_div_CryTmp_1_5_port, u_div_PartRem_1_1_port, 
      u_div_PartRem_1_2_port, u_div_PartRem_1_3_port, u_div_PartRem_1_4_port, 
      u_div_u_add_PartRem_3_0_SUM_4_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n7, Y => 
                           u_div_CryTmp_1_5_port);
   U2 : NOR2xp33_ASAP7_75t_R port map( A => n6, B => n10, Y => 
                           u_div_PartRem_1_4_port);
   U3 : INVx1_ASAP7_75t_R port map( A => a(0), Y => n1);
   U4 : NAND2xp33_ASAP7_75t_R port map( A => a(0), B => u_div_PartRem_1_1_port,
                           Y => n2);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n5, B => n2, Y => n3);
   U6 : OR2x2_ASAP7_75t_R port map( A => u_div_PartRem_1_3_port, B => n3, Y => 
                           n4);
   U7 : NOR2xp33_ASAP7_75t_R port map( A => n4, B => u_div_PartRem_1_4_port, Y 
                           => u_div_u_add_PartRem_3_0_SUM_4_port);
   U8 : XOR2xp5_ASAP7_75t_R port map( A => a(0), B => u_div_PartRem_1_1_port, Y
                           => u_div_SumTmp_0_1_port);
   U9 : XOR2xp5_ASAP7_75t_R port map( A => n5, B => n2, Y => 
                           u_div_SumTmp_0_2_port);
   U10 : XNOR2xp5_ASAP7_75t_R port map( A => u_div_PartRem_1_3_port, B => n3, Y
                           => u_div_SumTmp_0_3_port);
   U11 : XNOR2xp5_ASAP7_75t_R port map( A => u_div_PartRem_1_4_port, B => n4, Y
                           => u_div_SumTmp_0_4_port);
   U12 : INVx1_ASAP7_75t_R port map( A => u_div_PartRem_1_2_port, Y => n5);
   U13 : INVx1_ASAP7_75t_R port map( A => u_div_u_add_PartRem_3_0_SUM_4_port, Y
                           => u_div_CryTmp_0_6_port);
   U14 : INVx1_ASAP7_75t_R port map( A => n14, Y => u_div_MAdd_1_port);
   U15 : INVx1_ASAP7_75t_R port map( A => n13, Y => u_div_MAdd_2_port);
   U16 : INVx1_ASAP7_75t_R port map( A => n15, Y => u_div_MAdd_0_port);
   U17 : INVx1_ASAP7_75t_R port map( A => u_div_CryTmp_1_5_port, Y => n6);
   U18 : INVx1_ASAP7_75t_R port map( A => a(3), Y => n7);
   U19 : INVx1_ASAP7_75t_R port map( A => a(1), Y => n8);
   U20 : NAND3xp33_ASAP7_75t_R port map( A => n12, B => n17, C => n11, Y => n16
                           );
   U21 : NAND2xp33_ASAP7_75t_R port map( A => a(1), B => a(2), Y => n9);
   U22 : XOR2xp5_ASAP7_75t_R port map( A => a(1), B => a(2), Y => 
                           u_div_SumTmp_1_1_port);
   U23 : XNOR2xp5_ASAP7_75t_R port map( A => a(3), B => n9, Y => 
                           u_div_SumTmp_1_2_port);
   U24 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n7, Y => n10);
   U25 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_2_port, B => n16, Y => 
                           remainder(2));
   U26 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_1_port, B => n16, Y => 
                           remainder(1));
   U27 : AND2x2_ASAP7_75t_R port map( A => u_div_MAdd_0_port, B => n16, Y => 
                           remainder(0));
   U28 : AND3x1_ASAP7_75t_R port map( A => n15, B => n13, C => n14, Y => n17);
   U29 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_1_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_1_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n14);
   U30 : OAI22xp33_ASAP7_75t_R port map( A1 => a(1), A2 => n6, B1 => 
                           u_div_CryTmp_1_5_port, B2 => n8, Y => 
                           u_div_PartRem_1_1_port);
   U31 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_2_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_2_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n13);
   U32 : AO22x1_ASAP7_75t_R port map( A1 => u_div_SumTmp_1_1_port, A2 => 
                           u_div_CryTmp_1_5_port, B1 => a(2), B2 => n6, Y => 
                           u_div_PartRem_1_2_port);
   U33 : AOI22xp33_ASAP7_75t_R port map( A1 => n1, A2 => u_div_CryTmp_0_6_port,
                           B1 => u_div_u_add_PartRem_3_0_SUM_4_port, B2 => a(0)
                           , Y => n15);
   U34 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_3_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_3_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n12);
   U35 : AO22x1_ASAP7_75t_R port map( A1 => u_div_SumTmp_1_2_port, A2 => 
                           u_div_CryTmp_1_5_port, B1 => a(3), B2 => n6, Y => 
                           u_div_PartRem_1_3_port);
   U36 : AOI22xp33_ASAP7_75t_R port map( A1 => u_div_SumTmp_0_4_port, A2 => 
                           u_div_CryTmp_0_6_port, B1 => u_div_PartRem_1_4_port,
                           B2 => u_div_u_add_PartRem_3_0_SUM_4_port, Y => n11);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity dxyu_routing_Xis1_Yis1_Zis1_6 is

   port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;  
         routing : out std_logic_vector (6 downto 0));

end dxyu_routing_Xis1_Yis1_Zis1_6;

architecture SYN_rtl of dxyu_routing_Xis1_Yis1_Zis1_6 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND2xp5_ASAP7_75t_R port map( A => enable, B => n6, Y => n9);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => n3, B => n1, Y => n10);
   U19 : AND2x2_ASAP7_75t_R port map( A => n12, B => enable, Y => routing(6));
   U20 : NAND3xp33_ASAP7_75t_R port map( A => n2, B => n10, C => address(2), Y 
                           => n11);
   U21 : NAND3xp33_ASAP7_75t_R port map( A => n3, B => n4, C => enable, Y => n8
                           );
   U3 : NOR2xp33_ASAP7_75t_R port map( A => n10, B => n9, Y => routing(4));
   U4 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n3, Y => routing(2));
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n11, B => n7, Y => routing(5));
   U6 : NOR3xp33_ASAP7_75t_R port map( A => n5, B => address(1), C => n11, Y =>
                           routing(0));
   U7 : NOR4xp25_ASAP7_75t_R port map( A => address(2), B => n12, C => n8, D =>
                           n1, Y => routing(3));
   U9 : NOR2xp33_ASAP7_75t_R port map( A => address(0), B => address(1), Y => 
                           n12);
   U10 : NOR4xp25_ASAP7_75t_R port map( A => address(5), B => n9, C => n1, D =>
                           n4, Y => routing(1));
   U12 : INVx1_ASAP7_75t_R port map( A => address(4), Y => n1);
   U13 : INVx1_ASAP7_75t_R port map( A => n8, Y => n2);
   U14 : INVx1_ASAP7_75t_R port map( A => address(5), Y => n3);
   U15 : INVx1_ASAP7_75t_R port map( A => address(3), Y => n4);
   U16 : INVx1_ASAP7_75t_R port map( A => address(0), Y => n5);
   U17 : INVx1_ASAP7_75t_R port map( A => n12, Y => n6);
   U18 : INVx1_ASAP7_75t_R port map( A => address(1), Y => n7);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity dxyu_routing_Xis1_Yis1_Zis1_5 is

   port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;  
         routing : out std_logic_vector (6 downto 0));

end dxyu_routing_Xis1_Yis1_Zis1_5;

architecture SYN_rtl of dxyu_routing_Xis1_Yis1_Zis1_5 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND2xp5_ASAP7_75t_R port map( A => enable, B => n6, Y => n9);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => n3, B => n1, Y => n10);
   U19 : AND2x2_ASAP7_75t_R port map( A => n12, B => enable, Y => routing(6));
   U20 : NAND3xp33_ASAP7_75t_R port map( A => n2, B => n10, C => address(2), Y 
                           => n11);
   U21 : NAND3xp33_ASAP7_75t_R port map( A => n3, B => n4, C => enable, Y => n8
                           );
   U3 : NOR2xp33_ASAP7_75t_R port map( A => n10, B => n9, Y => routing(4));
   U4 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n3, Y => routing(2));
   U5 : NOR3xp33_ASAP7_75t_R port map( A => n5, B => address(1), C => n11, Y =>
                           routing(0));
   U6 : NOR2xp33_ASAP7_75t_R port map( A => n11, B => n7, Y => routing(5));
   U7 : NOR4xp25_ASAP7_75t_R port map( A => address(5), B => n9, C => n1, D => 
                           n4, Y => routing(1));
   U9 : NOR2xp33_ASAP7_75t_R port map( A => address(0), B => address(1), Y => 
                           n12);
   U10 : NOR4xp25_ASAP7_75t_R port map( A => address(2), B => n12, C => n8, D 
                           => n1, Y => routing(3));
   U12 : INVx1_ASAP7_75t_R port map( A => address(4), Y => n1);
   U13 : INVx1_ASAP7_75t_R port map( A => n8, Y => n2);
   U14 : INVx1_ASAP7_75t_R port map( A => address(5), Y => n3);
   U15 : INVx1_ASAP7_75t_R port map( A => address(3), Y => n4);
   U16 : INVx1_ASAP7_75t_R port map( A => address(0), Y => n5);
   U17 : INVx1_ASAP7_75t_R port map( A => n12, Y => n6);
   U18 : INVx1_ASAP7_75t_R port map( A => address(1), Y => n7);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity dxyu_routing_Xis1_Yis1_Zis1_4 is

   port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;  
         routing : out std_logic_vector (6 downto 0));

end dxyu_routing_Xis1_Yis1_Zis1_4;

architecture SYN_rtl of dxyu_routing_Xis1_Yis1_Zis1_4 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND2xp5_ASAP7_75t_R port map( A => enable, B => n6, Y => n9);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => n3, B => n1, Y => n10);
   U19 : AND2x2_ASAP7_75t_R port map( A => n12, B => enable, Y => routing(6));
   U20 : NAND3xp33_ASAP7_75t_R port map( A => n2, B => n10, C => address(2), Y 
                           => n11);
   U21 : NAND3xp33_ASAP7_75t_R port map( A => n3, B => n4, C => enable, Y => n8
                           );
   U3 : NOR2xp33_ASAP7_75t_R port map( A => n10, B => n9, Y => routing(4));
   U4 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n3, Y => routing(2));
   U5 : NOR3xp33_ASAP7_75t_R port map( A => n5, B => address(1), C => n11, Y =>
                           routing(0));
   U6 : NOR4xp25_ASAP7_75t_R port map( A => address(5), B => n9, C => n1, D => 
                           n4, Y => routing(1));
   U7 : NOR2xp33_ASAP7_75t_R port map( A => address(0), B => address(1), Y => 
                           n12);
   U9 : NOR2xp33_ASAP7_75t_R port map( A => n11, B => n7, Y => routing(5));
   U10 : NOR4xp25_ASAP7_75t_R port map( A => address(2), B => n12, C => n8, D 
                           => n1, Y => routing(3));
   U12 : INVx1_ASAP7_75t_R port map( A => address(4), Y => n1);
   U13 : INVx1_ASAP7_75t_R port map( A => n8, Y => n2);
   U14 : INVx1_ASAP7_75t_R port map( A => address(5), Y => n3);
   U15 : INVx1_ASAP7_75t_R port map( A => address(3), Y => n4);
   U16 : INVx1_ASAP7_75t_R port map( A => address(0), Y => n5);
   U17 : INVx1_ASAP7_75t_R port map( A => n12, Y => n6);
   U18 : INVx1_ASAP7_75t_R port map( A => address(1), Y => n7);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity dxyu_routing_Xis1_Yis1_Zis1_3 is

   port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;  
         routing : out std_logic_vector (6 downto 0));

end dxyu_routing_Xis1_Yis1_Zis1_3;

architecture SYN_rtl of dxyu_routing_Xis1_Yis1_Zis1_3 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND2xp5_ASAP7_75t_R port map( A => enable, B => n6, Y => n9);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => n3, B => n1, Y => n10);
   U19 : AND2x2_ASAP7_75t_R port map( A => n12, B => enable, Y => routing(6));
   U20 : NAND3xp33_ASAP7_75t_R port map( A => n2, B => n10, C => address(2), Y 
                           => n11);
   U21 : NAND3xp33_ASAP7_75t_R port map( A => n3, B => n4, C => enable, Y => n8
                           );
   U3 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n3, Y => routing(2));
   U4 : NOR2xp33_ASAP7_75t_R port map( A => n10, B => n9, Y => routing(4));
   U5 : NOR4xp25_ASAP7_75t_R port map( A => address(2), B => n12, C => n8, D =>
                           n1, Y => routing(3));
   U6 : NOR3xp33_ASAP7_75t_R port map( A => n5, B => address(1), C => n11, Y =>
                           routing(0));
   U7 : NOR4xp25_ASAP7_75t_R port map( A => address(5), B => n9, C => n1, D => 
                           n4, Y => routing(1));
   U9 : NOR2xp33_ASAP7_75t_R port map( A => address(0), B => address(1), Y => 
                           n12);
   U10 : NOR2xp33_ASAP7_75t_R port map( A => n11, B => n7, Y => routing(5));
   U12 : INVx1_ASAP7_75t_R port map( A => address(4), Y => n1);
   U13 : INVx1_ASAP7_75t_R port map( A => n8, Y => n2);
   U14 : INVx1_ASAP7_75t_R port map( A => address(5), Y => n3);
   U15 : INVx1_ASAP7_75t_R port map( A => address(3), Y => n4);
   U16 : INVx1_ASAP7_75t_R port map( A => address(0), Y => n5);
   U17 : INVx1_ASAP7_75t_R port map( A => n12, Y => n6);
   U18 : INVx1_ASAP7_75t_R port map( A => address(1), Y => n7);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity dxyu_routing_Xis1_Yis1_Zis1_2 is

   port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;  
         routing : out std_logic_vector (6 downto 0));

end dxyu_routing_Xis1_Yis1_Zis1_2;

architecture SYN_rtl of dxyu_routing_Xis1_Yis1_Zis1_2 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND2xp5_ASAP7_75t_R port map( A => enable, B => n6, Y => n9);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => n3, B => n1, Y => n10);
   U19 : AND2x2_ASAP7_75t_R port map( A => n12, B => enable, Y => routing(6));
   U20 : NAND3xp33_ASAP7_75t_R port map( A => n2, B => n10, C => address(2), Y 
                           => n11);
   U21 : NAND3xp33_ASAP7_75t_R port map( A => n3, B => n4, C => enable, Y => n8
                           );
   U3 : NOR2xp33_ASAP7_75t_R port map( A => n10, B => n9, Y => routing(4));
   U4 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n3, Y => routing(2));
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n11, B => n7, Y => routing(5));
   U6 : NOR4xp25_ASAP7_75t_R port map( A => address(2), B => n12, C => n8, D =>
                           n1, Y => routing(3));
   U7 : NOR2xp33_ASAP7_75t_R port map( A => address(0), B => address(1), Y => 
                           n12);
   U9 : NOR3xp33_ASAP7_75t_R port map( A => n5, B => address(1), C => n11, Y =>
                           routing(0));
   U10 : NOR4xp25_ASAP7_75t_R port map( A => address(5), B => n9, C => n1, D =>
                           n4, Y => routing(1));
   U12 : INVx1_ASAP7_75t_R port map( A => address(4), Y => n1);
   U13 : INVx1_ASAP7_75t_R port map( A => n8, Y => n2);
   U14 : INVx1_ASAP7_75t_R port map( A => address(5), Y => n3);
   U15 : INVx1_ASAP7_75t_R port map( A => address(3), Y => n4);
   U16 : INVx1_ASAP7_75t_R port map( A => address(0), Y => n5);
   U17 : INVx1_ASAP7_75t_R port map( A => n12, Y => n6);
   U18 : INVx1_ASAP7_75t_R port map( A => address(1), Y => n7);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity dxyu_routing_Xis1_Yis1_Zis1_1 is

   port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;  
         routing : out std_logic_vector (6 downto 0));

end dxyu_routing_Xis1_Yis1_Zis1_1;

architecture SYN_rtl of dxyu_routing_Xis1_Yis1_Zis1_1 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND2xp5_ASAP7_75t_R port map( A => enable, B => n6, Y => n9);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => n3, B => n1, Y => n10);
   U19 : AND2x2_ASAP7_75t_R port map( A => n12, B => enable, Y => routing(6));
   U20 : NAND3xp33_ASAP7_75t_R port map( A => n2, B => n10, C => address(2), Y 
                           => n11);
   U21 : NAND3xp33_ASAP7_75t_R port map( A => n3, B => n4, C => enable, Y => n8
                           );
   U3 : NOR2xp33_ASAP7_75t_R port map( A => n10, B => n9, Y => routing(4));
   U4 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => n3, Y => routing(2));
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n11, B => n7, Y => routing(5));
   U6 : NOR3xp33_ASAP7_75t_R port map( A => n5, B => address(1), C => n11, Y =>
                           routing(0));
   U7 : NOR2xp33_ASAP7_75t_R port map( A => address(0), B => address(1), Y => 
                           n12);
   U9 : NOR4xp25_ASAP7_75t_R port map( A => address(5), B => n9, C => n1, D => 
                           n4, Y => routing(1));
   U10 : NOR4xp25_ASAP7_75t_R port map( A => address(2), B => n12, C => n8, D 
                           => n1, Y => routing(3));
   U12 : INVx1_ASAP7_75t_R port map( A => address(4), Y => n1);
   U13 : INVx1_ASAP7_75t_R port map( A => n8, Y => n2);
   U14 : INVx1_ASAP7_75t_R port map( A => address(5), Y => n3);
   U15 : INVx1_ASAP7_75t_R port map( A => address(3), Y => n4);
   U16 : INVx1_ASAP7_75t_R port map( A => address(0), Y => n5);
   U17 : INVx1_ASAP7_75t_R port map( A => n12, Y => n6);
   U18 : INVx1_ASAP7_75t_R port map( A => address(1), Y => n7);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT6_6 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (5 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (5 downto 0));

end rr_arbiter_no_delay_CNT6_6;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT6_6 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AO21x1_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI31xp33_ASAP7_75t_R
      port( A1, A2, A3, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OR3x1_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO32x1_ASAP7_75t_R
      port( A1, A2, A3, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_5_port, grant_4_port, grant_3_port, grant_2_port, grant_1_port,
      grant_0_port, pre_req_5_port, pre_req_4_port, pre_req_3_port, 
      pre_req_2_port, pre_req_1_port, pre_req_0_port, N2, N3, N4, N5, N6, 
      mask_pre_5_port, mask_pre_4_port, mask_pre_3_port, mask_pre_2_port, N20, 
      n1, n2_port, n3_port, n4_port, n5_port, n8, n9, n10, n11, n12, n13, n15, 
      n17, n19, n21, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
      n50, n51, n52, n53, n54, n55 : std_logic;

begin
   grant <= ( grant_5_port, grant_4_port, grant_3_port, grant_2_port, 
      grant_1_port, grant_0_port );
   
   U13 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(5), A3 => n5_port, 
                           B1 => n15, B2 => mask_pre_5_port, Y => grant_5_port)
                           ;
   U14 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(4), A3 => n10, B1 =>
                           n21, B2 => mask_pre_4_port, Y => grant_4_port);
   U15 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(3), A3 => n9, B1 => 
                           n17, B2 => mask_pre_3_port, Y => grant_3_port);
   U16 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(2), A3 => n19, B1 =>
                           n8, B2 => mask_pre_2_port, Y => grant_2_port);
   U20 : OR3x1_ASAP7_75t_R port map( A => mask_pre_3_port, B => mask_pre_5_port
                           , C => mask_pre_4_port, Y => n54);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_4_port, A2 => ack, B1 => 
                           grant_4_port, B2 => n46, Y => n53);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_3_port, A2 => ack, B1 => 
                           grant_3_port, B2 => n46, Y => n52);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_2_port, A2 => ack, B1 => 
                           grant_2_port, B2 => n46, Y => n51);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_5_port, A2 => ack, B1 => 
                           grant_5_port, B2 => n46, Y => n50);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n46, Y => n49);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n46, Y => n48);
   pre_req_reg_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_4_port);
   pre_req_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_2_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n48, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_0_port);
   pre_req_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n52, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_3_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n49, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_1_port);
   pre_req_reg_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n50, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_5_port);
   U4 : TIELOx1_ASAP7_75t_R port map( L => n23);
   U5 : AND2x2_ASAP7_75t_R port map( A => n42, B => n40, Y => n1);
   U11 : AND2x2_ASAP7_75t_R port map( A => n43, B => n1, Y => n2_port);
   U12 : AND2x2_ASAP7_75t_R port map( A => n44, B => n2_port, Y => n3_port);
   U17 : AND2x2_ASAP7_75t_R port map( A => n39, B => n3_port, Y => n4_port);
   U18 : XOR2xp5_ASAP7_75t_R port map( A => n45, B => n4_port, Y => n5_port);
   U19 : XOR2xp5_ASAP7_75t_R port map( A => n36, B => n37, Y => n8);
   U21 : XOR2xp5_ASAP7_75t_R port map( A => n44, B => n2_port, Y => n9);
   U22 : XOR2xp5_ASAP7_75t_R port map( A => n39, B => n3_port, Y => n10);
   U23 : AND2x2_ASAP7_75t_R port map( A => n36, B => n37, Y => n11);
   U24 : AND2x2_ASAP7_75t_R port map( A => n35, B => n11, Y => n12);
   U25 : AND2x2_ASAP7_75t_R port map( A => n34, B => n12, Y => n13);
   U26 : XOR2xp5_ASAP7_75t_R port map( A => n33, B => n13, Y => n15);
   U27 : XOR2xp5_ASAP7_75t_R port map( A => n35, B => n11, Y => n17);
   U28 : XOR2xp5_ASAP7_75t_R port map( A => n43, B => n1, Y => n19);
   U29 : XOR2xp5_ASAP7_75t_R port map( A => n34, B => n12, Y => n21);
   U30 : NOR2xp33_ASAP7_75t_R port map( A => n41, B => n40, Y => grant_0_port);
   U31 : NOR3xp33_ASAP7_75t_R port map( A => n54, B => N20, C => 
                           mask_pre_2_port, Y => n55);
   U32 : INVx1_ASAP7_75t_R port map( A => rst, Y => n25);
   U33 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_2_port, B => N3, C => n43,
                           Y => mask_pre_2_port);
   U34 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_1_port, B => N2, C => n42,
                           Y => N20);
   U35 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_3_port, B => N4, C => n44,
                           Y => mask_pre_3_port);
   U36 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_5_port, B => N6, C => n45,
                           Y => mask_pre_5_port);
   U37 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_4_port, B => N5, C => n47,
                           Y => mask_pre_4_port);
   U38 : OAI31xp33_ASAP7_75t_R port map( A1 => n41, A2 => n38, A3 => n42, B => 
                           n37, Y => grant_1_port);
   U39 : XNOR2xp5_ASAP7_75t_R port map( A => n42, B => n40, Y => n38);
   U40 : NOR2xp33_ASAP7_75t_R port map( A => pre_req_1_port, B => 
                           pre_req_0_port, Y => n26);
   U41 : AO21x1_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => 
                           pre_req_1_port, B => n26, Y => N2);
   U42 : NOR2xp33_ASAP7_75t_R port map( A => n30, B => pre_req_2_port, Y => n27
                           );
   U43 : AO21x1_ASAP7_75t_R port map( A1 => n30, A2 => pre_req_2_port, B => n27
                           , Y => N3);
   U44 : NOR2xp33_ASAP7_75t_R port map( A => n31, B => pre_req_3_port, Y => n28
                           );
   U45 : AO21x1_ASAP7_75t_R port map( A1 => n31, A2 => pre_req_3_port, B => n28
                           , Y => N4);
   U46 : XNOR2xp5_ASAP7_75t_R port map( A => pre_req_4_port, B => n32, Y => N5)
                           ;
   U47 : NOR2xp33_ASAP7_75t_R port map( A => pre_req_4_port, B => n32, Y => n29
                           );
   U48 : XOR2xp5_ASAP7_75t_R port map( A => pre_req_5_port, B => n29, Y => N6);
   U49 : INVx1_ASAP7_75t_R port map( A => n26, Y => n30);
   U50 : INVx1_ASAP7_75t_R port map( A => n27, Y => n31);
   U51 : INVx1_ASAP7_75t_R port map( A => n28, Y => n32);
   U52 : INVx1_ASAP7_75t_R port map( A => mask_pre_5_port, Y => n33);
   U53 : INVx1_ASAP7_75t_R port map( A => mask_pre_4_port, Y => n34);
   U54 : INVx1_ASAP7_75t_R port map( A => mask_pre_3_port, Y => n35);
   U55 : INVx1_ASAP7_75t_R port map( A => mask_pre_2_port, Y => n36);
   U56 : INVx1_ASAP7_75t_R port map( A => N20, Y => n37);
   U57 : INVx1_ASAP7_75t_R port map( A => req(4), Y => n39);
   U58 : INVx1_ASAP7_75t_R port map( A => req(0), Y => n40);
   U59 : INVx1_ASAP7_75t_R port map( A => n55, Y => n41);
   U60 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n42);
   U61 : INVx1_ASAP7_75t_R port map( A => req(2), Y => n43);
   U62 : INVx1_ASAP7_75t_R port map( A => req(3), Y => n44);
   U63 : INVx1_ASAP7_75t_R port map( A => req(5), Y => n45);
   U64 : INVx1_ASAP7_75t_R port map( A => ack, Y => n46);
   U65 : INVx1_ASAP7_75t_R port map( A => req(4), Y => n47);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT6_5 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (5 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (5 downto 0));

end rr_arbiter_no_delay_CNT6_5;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT6_5 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AO21x1_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI31xp33_ASAP7_75t_R
      port( A1, A2, A3, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OR3x1_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO32x1_ASAP7_75t_R
      port( A1, A2, A3, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_5_port, grant_4_port, grant_3_port, grant_2_port, grant_1_port,
      grant_0_port, pre_req_5_port, pre_req_4_port, pre_req_3_port, 
      pre_req_2_port, pre_req_1_port, pre_req_0_port, N2, N3, N4, N5, N6, 
      mask_pre_5_port, mask_pre_4_port, mask_pre_3_port, mask_pre_2_port, N20, 
      n1, n2_port, n3_port, n4_port, n5_port, n8, n9, n10, n11, n12, n13, n15, 
      n17, n19, n21, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
      n50, n51, n52, n53, n54, n55, n56 : std_logic;

begin
   grant <= ( grant_5_port, grant_4_port, grant_3_port, grant_2_port, 
      grant_1_port, grant_0_port );
   
   U13 : AO32x1_ASAP7_75t_R port map( A1 => n56, A2 => req(5), A3 => n9, B1 => 
                           n21, B2 => mask_pre_5_port, Y => grant_5_port);
   U14 : AO32x1_ASAP7_75t_R port map( A1 => n56, A2 => req(4), A3 => n4_port, 
                           B1 => n12, B2 => mask_pre_4_port, Y => grant_4_port)
                           ;
   U15 : AO32x1_ASAP7_75t_R port map( A1 => n56, A2 => req(3), A3 => n8, B1 => 
                           n19, B2 => mask_pre_3_port, Y => grant_3_port);
   U16 : AO32x1_ASAP7_75t_R port map( A1 => n56, A2 => req(2), A3 => n13, B1 =>
                           n5_port, B2 => mask_pre_2_port, Y => grant_2_port);
   U20 : OR3x1_ASAP7_75t_R port map( A => mask_pre_3_port, B => mask_pre_5_port
                           , C => mask_pre_4_port, Y => n55);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_4_port, A2 => ack, B1 => 
                           grant_4_port, B2 => n45, Y => n54);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_3_port, A2 => ack, B1 => 
                           grant_3_port, B2 => n45, Y => n53);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_2_port, A2 => ack, B1 => 
                           grant_2_port, B2 => n45, Y => n52);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_5_port, A2 => ack, B1 => 
                           grant_5_port, B2 => n45, Y => n51);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n45, Y => n50);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n45, Y => n49);
   pre_req_reg_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_5_port);
   pre_req_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_3_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n49, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_0_port);
   pre_req_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n52, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_2_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n50, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_1_port);
   pre_req_reg_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n54, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_4_port);
   U4 : TIELOx1_ASAP7_75t_R port map( L => n23);
   U5 : AND2x2_ASAP7_75t_R port map( A => n40, B => n3_port, Y => n1);
   U11 : AND2x2_ASAP7_75t_R port map( A => n42, B => n41, Y => n2_port);
   U12 : AND2x2_ASAP7_75t_R port map( A => n44, B => n2_port, Y => n3_port);
   U17 : XOR2xp5_ASAP7_75t_R port map( A => n46, B => n1, Y => n4_port);
   U18 : XOR2xp5_ASAP7_75t_R port map( A => n36, B => n37, Y => n5_port);
   U19 : XOR2xp5_ASAP7_75t_R port map( A => n40, B => n3_port, Y => n8);
   U21 : XOR2xp5_ASAP7_75t_R port map( A => n39, B => n17, Y => n9);
   U22 : AND2x2_ASAP7_75t_R port map( A => n36, B => n37, Y => n10);
   U23 : AND2x2_ASAP7_75t_R port map( A => n35, B => n10, Y => n11);
   U24 : XOR2xp5_ASAP7_75t_R port map( A => n34, B => n11, Y => n12);
   U25 : XOR2xp5_ASAP7_75t_R port map( A => n44, B => n2_port, Y => n13);
   U26 : AND2x2_ASAP7_75t_R port map( A => n34, B => n11, Y => n15);
   U27 : AND2x2_ASAP7_75t_R port map( A => n46, B => n1, Y => n17);
   U28 : XOR2xp5_ASAP7_75t_R port map( A => n35, B => n10, Y => n19);
   U29 : XOR2xp5_ASAP7_75t_R port map( A => n33, B => n15, Y => n21);
   U30 : NOR3xp33_ASAP7_75t_R port map( A => n55, B => N20, C => 
                           mask_pre_2_port, Y => n56);
   U31 : INVx1_ASAP7_75t_R port map( A => rst, Y => n25);
   U32 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_2_port, B => N3, C => n44,
                           Y => mask_pre_2_port);
   U33 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_1_port, B => N2, C => n42,
                           Y => N20);
   U34 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_4_port, B => N5, C => n46,
                           Y => mask_pre_4_port);
   U35 : NOR2xp33_ASAP7_75t_R port map( A => n43, B => n41, Y => grant_0_port);
   U36 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_5_port, B => N6, C => n48,
                           Y => mask_pre_5_port);
   U37 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_3_port, B => N4, C => n47,
                           Y => mask_pre_3_port);
   U38 : OAI31xp33_ASAP7_75t_R port map( A1 => n43, A2 => n38, A3 => n42, B => 
                           n37, Y => grant_1_port);
   U39 : XNOR2xp5_ASAP7_75t_R port map( A => n42, B => n41, Y => n38);
   U40 : NOR2xp33_ASAP7_75t_R port map( A => pre_req_1_port, B => 
                           pre_req_0_port, Y => n26);
   U41 : AO21x1_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => 
                           pre_req_1_port, B => n26, Y => N2);
   U42 : NOR2xp33_ASAP7_75t_R port map( A => n30, B => pre_req_2_port, Y => n27
                           );
   U43 : AO21x1_ASAP7_75t_R port map( A1 => n30, A2 => pre_req_2_port, B => n27
                           , Y => N3);
   U44 : NOR2xp33_ASAP7_75t_R port map( A => n31, B => pre_req_3_port, Y => n28
                           );
   U45 : AO21x1_ASAP7_75t_R port map( A1 => n31, A2 => pre_req_3_port, B => n28
                           , Y => N4);
   U46 : XNOR2xp5_ASAP7_75t_R port map( A => pre_req_4_port, B => n32, Y => N5)
                           ;
   U47 : NOR2xp33_ASAP7_75t_R port map( A => pre_req_4_port, B => n32, Y => n29
                           );
   U48 : XOR2xp5_ASAP7_75t_R port map( A => pre_req_5_port, B => n29, Y => N6);
   U49 : INVx1_ASAP7_75t_R port map( A => n26, Y => n30);
   U50 : INVx1_ASAP7_75t_R port map( A => n27, Y => n31);
   U51 : INVx1_ASAP7_75t_R port map( A => n28, Y => n32);
   U52 : INVx1_ASAP7_75t_R port map( A => mask_pre_5_port, Y => n33);
   U53 : INVx1_ASAP7_75t_R port map( A => mask_pre_4_port, Y => n34);
   U54 : INVx1_ASAP7_75t_R port map( A => mask_pre_3_port, Y => n35);
   U55 : INVx1_ASAP7_75t_R port map( A => mask_pre_2_port, Y => n36);
   U56 : INVx1_ASAP7_75t_R port map( A => N20, Y => n37);
   U57 : INVx1_ASAP7_75t_R port map( A => req(5), Y => n39);
   U58 : INVx1_ASAP7_75t_R port map( A => req(3), Y => n40);
   U59 : INVx1_ASAP7_75t_R port map( A => req(0), Y => n41);
   U60 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n42);
   U61 : INVx1_ASAP7_75t_R port map( A => n56, Y => n43);
   U62 : INVx1_ASAP7_75t_R port map( A => req(2), Y => n44);
   U63 : INVx1_ASAP7_75t_R port map( A => ack, Y => n45);
   U64 : INVx1_ASAP7_75t_R port map( A => req(4), Y => n46);
   U65 : INVx1_ASAP7_75t_R port map( A => req(3), Y => n47);
   U66 : INVx1_ASAP7_75t_R port map( A => req(5), Y => n48);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT6_4 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (5 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (5 downto 0));

end rr_arbiter_no_delay_CNT6_4;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT6_4 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AO21x1_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI31xp33_ASAP7_75t_R
      port( A1, A2, A3, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OR3x1_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO32x1_ASAP7_75t_R
      port( A1, A2, A3, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_5_port, grant_4_port, grant_3_port, grant_2_port, grant_1_port,
      grant_0_port, pre_req_5_port, pre_req_4_port, pre_req_3_port, 
      pre_req_2_port, pre_req_1_port, pre_req_0_port, N2, N3, N4, N5, N6, 
      mask_pre_5_port, mask_pre_4_port, mask_pre_3_port, mask_pre_2_port, N20, 
      n1, n2_port, n3_port, n4_port, n5_port, n8, n9, n10, n11, n12, n13, n15, 
      n17, n19, n21, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
      n50, n51, n52, n53, n54, n55 : std_logic;

begin
   grant <= ( grant_5_port, grant_4_port, grant_3_port, grant_2_port, 
      grant_1_port, grant_0_port );
   
   U13 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(5), A3 => n4_port, 
                           B1 => n13, B2 => mask_pre_5_port, Y => grant_5_port)
                           ;
   U14 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(4), A3 => n5_port, 
                           B1 => n17, B2 => mask_pre_4_port, Y => grant_4_port)
                           ;
   U15 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(3), A3 => n8, B1 => 
                           n19, B2 => mask_pre_3_port, Y => grant_3_port);
   U16 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(2), A3 => n9, B1 => 
                           n21, B2 => mask_pre_2_port, Y => grant_2_port);
   U20 : OR3x1_ASAP7_75t_R port map( A => mask_pre_3_port, B => mask_pre_5_port
                           , C => mask_pre_4_port, Y => n54);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_4_port, A2 => ack, B1 => 
                           grant_4_port, B2 => n45, Y => n53);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_3_port, A2 => ack, B1 => 
                           grant_3_port, B2 => n45, Y => n52);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_2_port, A2 => ack, B1 => 
                           grant_2_port, B2 => n45, Y => n51);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_5_port, A2 => ack, B1 => 
                           grant_5_port, B2 => n45, Y => n50);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n45, Y => n49);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n45, Y => n48);
   pre_req_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_2_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n49, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n48, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_0_port);
   pre_req_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n52, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_3_port);
   pre_req_reg_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_4_port);
   pre_req_reg_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n50, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_5_port);
   U4 : TIELOx1_ASAP7_75t_R port map( L => n23);
   U5 : AND2x2_ASAP7_75t_R port map( A => n46, B => n2_port, Y => n1);
   U11 : AND2x2_ASAP7_75t_R port map( A => n39, B => n15, Y => n2_port);
   U12 : AND2x2_ASAP7_75t_R port map( A => n42, B => n1, Y => n3_port);
   U17 : XOR2xp5_ASAP7_75t_R port map( A => n43, B => n3_port, Y => n4_port);
   U18 : XOR2xp5_ASAP7_75t_R port map( A => n42, B => n1, Y => n5_port);
   U19 : XOR2xp5_ASAP7_75t_R port map( A => n46, B => n2_port, Y => n8);
   U21 : XOR2xp5_ASAP7_75t_R port map( A => n39, B => n15, Y => n9);
   U22 : AND2x2_ASAP7_75t_R port map( A => n36, B => n37, Y => n10);
   U23 : AND2x2_ASAP7_75t_R port map( A => n35, B => n10, Y => n11);
   U24 : AND2x2_ASAP7_75t_R port map( A => n34, B => n11, Y => n12);
   U25 : XOR2xp5_ASAP7_75t_R port map( A => n33, B => n12, Y => n13);
   U26 : AND2x2_ASAP7_75t_R port map( A => n44, B => n40, Y => n15);
   U27 : XOR2xp5_ASAP7_75t_R port map( A => n34, B => n11, Y => n17);
   U28 : XOR2xp5_ASAP7_75t_R port map( A => n35, B => n10, Y => n19);
   U29 : XOR2xp5_ASAP7_75t_R port map( A => n36, B => n37, Y => n21);
   U30 : NOR2xp33_ASAP7_75t_R port map( A => n41, B => n40, Y => grant_0_port);
   U31 : NOR3xp33_ASAP7_75t_R port map( A => n54, B => N20, C => 
                           mask_pre_2_port, Y => n55);
   U32 : INVx1_ASAP7_75t_R port map( A => rst, Y => n25);
   U33 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_1_port, B => N2, C => n44,
                           Y => N20);
   U34 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_5_port, B => N6, C => n43,
                           Y => mask_pre_5_port);
   U35 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_4_port, B => N5, C => n42,
                           Y => mask_pre_4_port);
   U36 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_3_port, B => N4, C => n46,
                           Y => mask_pre_3_port);
   U37 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_2_port, B => N3, C => n47,
                           Y => mask_pre_2_port);
   U38 : OAI31xp33_ASAP7_75t_R port map( A1 => n41, A2 => n38, A3 => n44, B => 
                           n37, Y => grant_1_port);
   U39 : XNOR2xp5_ASAP7_75t_R port map( A => n44, B => n40, Y => n38);
   U40 : NOR2xp33_ASAP7_75t_R port map( A => pre_req_1_port, B => 
                           pre_req_0_port, Y => n26);
   U41 : AO21x1_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => 
                           pre_req_1_port, B => n26, Y => N2);
   U42 : NOR2xp33_ASAP7_75t_R port map( A => n30, B => pre_req_2_port, Y => n27
                           );
   U43 : AO21x1_ASAP7_75t_R port map( A1 => n30, A2 => pre_req_2_port, B => n27
                           , Y => N3);
   U44 : NOR2xp33_ASAP7_75t_R port map( A => n31, B => pre_req_3_port, Y => n28
                           );
   U45 : AO21x1_ASAP7_75t_R port map( A1 => n31, A2 => pre_req_3_port, B => n28
                           , Y => N4);
   U46 : XNOR2xp5_ASAP7_75t_R port map( A => pre_req_4_port, B => n32, Y => N5)
                           ;
   U47 : NOR2xp33_ASAP7_75t_R port map( A => pre_req_4_port, B => n32, Y => n29
                           );
   U48 : XOR2xp5_ASAP7_75t_R port map( A => pre_req_5_port, B => n29, Y => N6);
   U49 : INVx1_ASAP7_75t_R port map( A => n26, Y => n30);
   U50 : INVx1_ASAP7_75t_R port map( A => n27, Y => n31);
   U51 : INVx1_ASAP7_75t_R port map( A => n28, Y => n32);
   U52 : INVx1_ASAP7_75t_R port map( A => mask_pre_5_port, Y => n33);
   U53 : INVx1_ASAP7_75t_R port map( A => mask_pre_4_port, Y => n34);
   U54 : INVx1_ASAP7_75t_R port map( A => mask_pre_3_port, Y => n35);
   U55 : INVx1_ASAP7_75t_R port map( A => mask_pre_2_port, Y => n36);
   U56 : INVx1_ASAP7_75t_R port map( A => N20, Y => n37);
   U57 : INVx1_ASAP7_75t_R port map( A => req(2), Y => n39);
   U58 : INVx1_ASAP7_75t_R port map( A => req(0), Y => n40);
   U59 : INVx1_ASAP7_75t_R port map( A => n55, Y => n41);
   U60 : INVx1_ASAP7_75t_R port map( A => req(4), Y => n42);
   U61 : INVx1_ASAP7_75t_R port map( A => req(5), Y => n43);
   U62 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n44);
   U63 : INVx1_ASAP7_75t_R port map( A => ack, Y => n45);
   U64 : INVx1_ASAP7_75t_R port map( A => req(3), Y => n46);
   U65 : INVx1_ASAP7_75t_R port map( A => req(2), Y => n47);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT6_3 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (5 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (5 downto 0));

end rr_arbiter_no_delay_CNT6_3;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT6_3 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AO21x1_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI31xp33_ASAP7_75t_R
      port( A1, A2, A3, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OR3x1_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO32x1_ASAP7_75t_R
      port( A1, A2, A3, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_5_port, grant_4_port, grant_3_port, grant_2_port, grant_1_port,
      grant_0_port, pre_req_5_port, pre_req_4_port, pre_req_3_port, 
      pre_req_2_port, pre_req_1_port, pre_req_0_port, N2, N3, N4, N5, N6, 
      mask_pre_5_port, mask_pre_4_port, mask_pre_3_port, mask_pre_2_port, N20, 
      n1, n2_port, n3_port, n4_port, n5_port, n8, n9, n10, n11, n12, n13, n15, 
      n17, n19, n21, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
      n50, n51, n52, n53, n54, n55 : std_logic;

begin
   grant <= ( grant_5_port, grant_4_port, grant_3_port, grant_2_port, 
      grant_1_port, grant_0_port );
   
   U13 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(5), A3 => n10, B1 =>
                           n21, B2 => mask_pre_5_port, Y => grant_5_port);
   U14 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(4), A3 => n4_port, 
                           B1 => n11, B2 => mask_pre_4_port, Y => grant_4_port)
                           ;
   U15 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(3), A3 => n9, B1 => 
                           n19, B2 => mask_pre_3_port, Y => grant_3_port);
   U16 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(2), A3 => n5_port, 
                           B1 => n13, B2 => mask_pre_2_port, Y => grant_2_port)
                           ;
   U20 : OR3x1_ASAP7_75t_R port map( A => mask_pre_3_port, B => mask_pre_5_port
                           , C => mask_pre_4_port, Y => n54);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_4_port, A2 => ack, B1 => 
                           grant_4_port, B2 => n45, Y => n53);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_3_port, A2 => ack, B1 => 
                           grant_3_port, B2 => n45, Y => n52);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_2_port, A2 => ack, B1 => 
                           grant_2_port, B2 => n45, Y => n51);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_5_port, A2 => ack, B1 => 
                           grant_5_port, B2 => n45, Y => n50);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n45, Y => n49);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n45, Y => n48);
   pre_req_reg_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n50, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_5_port);
   pre_req_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n52, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_3_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n49, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_1_port);
   pre_req_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_2_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n48, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_0_port);
   pre_req_reg_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_4_port);
   U4 : TIELOx1_ASAP7_75t_R port map( L => n23);
   U5 : AND2x2_ASAP7_75t_R port map( A => n40, B => n3_port, Y => n1);
   U11 : AND2x2_ASAP7_75t_R port map( A => n41, B => n42, Y => n2_port);
   U12 : AND2x2_ASAP7_75t_R port map( A => n46, B => n2_port, Y => n3_port);
   U17 : XOR2xp5_ASAP7_75t_R port map( A => n44, B => n1, Y => n4_port);
   U18 : XOR2xp5_ASAP7_75t_R port map( A => n46, B => n2_port, Y => n5_port);
   U19 : AND2x2_ASAP7_75t_R port map( A => n35, B => n12, Y => n8);
   U21 : XOR2xp5_ASAP7_75t_R port map( A => n40, B => n3_port, Y => n9);
   U22 : XOR2xp5_ASAP7_75t_R port map( A => n39, B => n17, Y => n10);
   U23 : XOR2xp5_ASAP7_75t_R port map( A => n34, B => n8, Y => n11);
   U24 : AND2x2_ASAP7_75t_R port map( A => n36, B => n37, Y => n12);
   U25 : XOR2xp5_ASAP7_75t_R port map( A => n36, B => n37, Y => n13);
   U26 : AND2x2_ASAP7_75t_R port map( A => n34, B => n8, Y => n15);
   U27 : AND2x2_ASAP7_75t_R port map( A => n44, B => n1, Y => n17);
   U28 : XOR2xp5_ASAP7_75t_R port map( A => n35, B => n12, Y => n19);
   U29 : XOR2xp5_ASAP7_75t_R port map( A => n33, B => n15, Y => n21);
   U30 : NOR2xp33_ASAP7_75t_R port map( A => n43, B => n42, Y => grant_0_port);
   U31 : NOR3xp33_ASAP7_75t_R port map( A => n54, B => N20, C => 
                           mask_pre_2_port, Y => n55);
   U32 : INVx1_ASAP7_75t_R port map( A => rst, Y => n25);
   U33 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_4_port, B => N5, C => n44,
                           Y => mask_pre_4_port);
   U34 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_2_port, B => N3, C => n46,
                           Y => mask_pre_2_port);
   U35 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_1_port, B => N2, C => n47,
                           Y => N20);
   U36 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_5_port, B => N6, C => n39,
                           Y => mask_pre_5_port);
   U37 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_3_port, B => N4, C => n40,
                           Y => mask_pre_3_port);
   U38 : OAI31xp33_ASAP7_75t_R port map( A1 => n43, A2 => n38, A3 => n47, B => 
                           n37, Y => grant_1_port);
   U39 : XNOR2xp5_ASAP7_75t_R port map( A => n41, B => n42, Y => n38);
   U40 : NOR2xp33_ASAP7_75t_R port map( A => pre_req_1_port, B => 
                           pre_req_0_port, Y => n26);
   U41 : AO21x1_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => 
                           pre_req_1_port, B => n26, Y => N2);
   U42 : NOR2xp33_ASAP7_75t_R port map( A => n30, B => pre_req_2_port, Y => n27
                           );
   U43 : AO21x1_ASAP7_75t_R port map( A1 => n30, A2 => pre_req_2_port, B => n27
                           , Y => N3);
   U44 : NOR2xp33_ASAP7_75t_R port map( A => n31, B => pre_req_3_port, Y => n28
                           );
   U45 : AO21x1_ASAP7_75t_R port map( A1 => n31, A2 => pre_req_3_port, B => n28
                           , Y => N4);
   U46 : XNOR2xp5_ASAP7_75t_R port map( A => pre_req_4_port, B => n32, Y => N5)
                           ;
   U47 : NOR2xp33_ASAP7_75t_R port map( A => pre_req_4_port, B => n32, Y => n29
                           );
   U48 : XOR2xp5_ASAP7_75t_R port map( A => pre_req_5_port, B => n29, Y => N6);
   U49 : INVx1_ASAP7_75t_R port map( A => n26, Y => n30);
   U50 : INVx1_ASAP7_75t_R port map( A => n27, Y => n31);
   U51 : INVx1_ASAP7_75t_R port map( A => n28, Y => n32);
   U52 : INVx1_ASAP7_75t_R port map( A => mask_pre_5_port, Y => n33);
   U53 : INVx1_ASAP7_75t_R port map( A => mask_pre_4_port, Y => n34);
   U54 : INVx1_ASAP7_75t_R port map( A => mask_pre_3_port, Y => n35);
   U55 : INVx1_ASAP7_75t_R port map( A => mask_pre_2_port, Y => n36);
   U56 : INVx1_ASAP7_75t_R port map( A => N20, Y => n37);
   U57 : INVx1_ASAP7_75t_R port map( A => req(5), Y => n39);
   U58 : INVx1_ASAP7_75t_R port map( A => req(3), Y => n40);
   U59 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n41);
   U60 : INVx1_ASAP7_75t_R port map( A => req(0), Y => n42);
   U61 : INVx1_ASAP7_75t_R port map( A => n55, Y => n43);
   U62 : INVx1_ASAP7_75t_R port map( A => req(4), Y => n44);
   U63 : INVx1_ASAP7_75t_R port map( A => ack, Y => n45);
   U64 : INVx1_ASAP7_75t_R port map( A => req(2), Y => n46);
   U65 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n47);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT6_2 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (5 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (5 downto 0));

end rr_arbiter_no_delay_CNT6_2;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT6_2 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AO21x1_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI31xp33_ASAP7_75t_R
      port( A1, A2, A3, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OR3x1_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO32x1_ASAP7_75t_R
      port( A1, A2, A3, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_5_port, grant_4_port, grant_3_port, grant_2_port, grant_1_port,
      grant_0_port, pre_req_5_port, pre_req_4_port, pre_req_3_port, 
      pre_req_2_port, pre_req_1_port, pre_req_0_port, N2, N3, N4, N5, N6, 
      mask_pre_5_port, mask_pre_4_port, mask_pre_3_port, mask_pre_2_port, N20, 
      n1, n2_port, n3_port, n4_port, n5_port, n8, n9, n10, n11, n12, n13, n15, 
      n17, n19, n21, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
      n50, n51, n52, n53, n54 : std_logic;

begin
   grant <= ( grant_5_port, grant_4_port, grant_3_port, grant_2_port, 
      grant_1_port, grant_0_port );
   
   U13 : AO32x1_ASAP7_75t_R port map( A1 => n54, A2 => req(5), A3 => n5_port, 
                           B1 => n15, B2 => mask_pre_5_port, Y => grant_5_port)
                           ;
   U14 : AO32x1_ASAP7_75t_R port map( A1 => n54, A2 => req(4), A3 => n9, B1 => 
                           n17, B2 => mask_pre_4_port, Y => grant_4_port);
   U15 : AO32x1_ASAP7_75t_R port map( A1 => n54, A2 => req(3), A3 => n19, B1 =>
                           n8, B2 => mask_pre_3_port, Y => grant_3_port);
   U16 : AO32x1_ASAP7_75t_R port map( A1 => n54, A2 => req(2), A3 => n21, B1 =>
                           n10, B2 => mask_pre_2_port, Y => grant_2_port);
   U20 : OR3x1_ASAP7_75t_R port map( A => mask_pre_3_port, B => mask_pre_5_port
                           , C => mask_pre_4_port, Y => n53);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_4_port, A2 => ack, B1 => 
                           grant_4_port, B2 => n45, Y => n52);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_3_port, A2 => ack, B1 => 
                           grant_3_port, B2 => n45, Y => n51);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_2_port, A2 => ack, B1 => 
                           grant_2_port, B2 => n45, Y => n50);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_5_port, A2 => ack, B1 => 
                           grant_5_port, B2 => n45, Y => n49);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n45, Y => n48);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n45, Y => n47);
   pre_req_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n50, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_2_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n48, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n47, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_0_port);
   pre_req_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_3_port);
   pre_req_reg_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n52, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_4_port);
   pre_req_reg_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n49, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_5_port);
   U4 : TIELOx1_ASAP7_75t_R port map( L => n23);
   U5 : AND2x2_ASAP7_75t_R port map( A => n46, B => n39, Y => n1);
   U11 : AND2x2_ASAP7_75t_R port map( A => n41, B => n1, Y => n2_port);
   U12 : AND2x2_ASAP7_75t_R port map( A => n42, B => n2_port, Y => n3_port);
   U17 : AND2x2_ASAP7_75t_R port map( A => n43, B => n3_port, Y => n4_port);
   U18 : XOR2xp5_ASAP7_75t_R port map( A => n44, B => n4_port, Y => n5_port);
   U19 : XOR2xp5_ASAP7_75t_R port map( A => n35, B => n11, Y => n8);
   U21 : XOR2xp5_ASAP7_75t_R port map( A => n43, B => n3_port, Y => n9);
   U22 : XOR2xp5_ASAP7_75t_R port map( A => n36, B => n37, Y => n10);
   U23 : AND2x2_ASAP7_75t_R port map( A => n36, B => n37, Y => n11);
   U24 : AND2x2_ASAP7_75t_R port map( A => n35, B => n11, Y => n12);
   U25 : AND2x2_ASAP7_75t_R port map( A => n34, B => n12, Y => n13);
   U26 : XOR2xp5_ASAP7_75t_R port map( A => n33, B => n13, Y => n15);
   U27 : XOR2xp5_ASAP7_75t_R port map( A => n34, B => n12, Y => n17);
   U28 : XOR2xp5_ASAP7_75t_R port map( A => n42, B => n2_port, Y => n19);
   U29 : XOR2xp5_ASAP7_75t_R port map( A => n41, B => n1, Y => n21);
   U30 : NOR2xp33_ASAP7_75t_R port map( A => n40, B => n39, Y => grant_0_port);
   U31 : NOR3xp33_ASAP7_75t_R port map( A => n53, B => N20, C => 
                           mask_pre_2_port, Y => n54);
   U32 : INVx1_ASAP7_75t_R port map( A => rst, Y => n25);
   U33 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_2_port, B => N3, C => n41,
                           Y => mask_pre_2_port);
   U34 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_3_port, B => N4, C => n42,
                           Y => mask_pre_3_port);
   U35 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_4_port, B => N5, C => n43,
                           Y => mask_pre_4_port);
   U36 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_5_port, B => N6, C => n44,
                           Y => mask_pre_5_port);
   U37 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_1_port, B => N2, C => n46,
                           Y => N20);
   U38 : OAI31xp33_ASAP7_75t_R port map( A1 => n40, A2 => n38, A3 => n46, B => 
                           n37, Y => grant_1_port);
   U39 : XNOR2xp5_ASAP7_75t_R port map( A => n46, B => n39, Y => n38);
   U40 : NOR2xp33_ASAP7_75t_R port map( A => pre_req_1_port, B => 
                           pre_req_0_port, Y => n26);
   U41 : AO21x1_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => 
                           pre_req_1_port, B => n26, Y => N2);
   U42 : NOR2xp33_ASAP7_75t_R port map( A => n30, B => pre_req_2_port, Y => n27
                           );
   U43 : AO21x1_ASAP7_75t_R port map( A1 => n30, A2 => pre_req_2_port, B => n27
                           , Y => N3);
   U44 : NOR2xp33_ASAP7_75t_R port map( A => n31, B => pre_req_3_port, Y => n28
                           );
   U45 : AO21x1_ASAP7_75t_R port map( A1 => n31, A2 => pre_req_3_port, B => n28
                           , Y => N4);
   U46 : XNOR2xp5_ASAP7_75t_R port map( A => pre_req_4_port, B => n32, Y => N5)
                           ;
   U47 : NOR2xp33_ASAP7_75t_R port map( A => pre_req_4_port, B => n32, Y => n29
                           );
   U48 : XOR2xp5_ASAP7_75t_R port map( A => pre_req_5_port, B => n29, Y => N6);
   U49 : INVx1_ASAP7_75t_R port map( A => n26, Y => n30);
   U50 : INVx1_ASAP7_75t_R port map( A => n27, Y => n31);
   U51 : INVx1_ASAP7_75t_R port map( A => n28, Y => n32);
   U52 : INVx1_ASAP7_75t_R port map( A => mask_pre_5_port, Y => n33);
   U53 : INVx1_ASAP7_75t_R port map( A => mask_pre_4_port, Y => n34);
   U54 : INVx1_ASAP7_75t_R port map( A => mask_pre_3_port, Y => n35);
   U55 : INVx1_ASAP7_75t_R port map( A => mask_pre_2_port, Y => n36);
   U56 : INVx1_ASAP7_75t_R port map( A => N20, Y => n37);
   U57 : INVx1_ASAP7_75t_R port map( A => req(0), Y => n39);
   U58 : INVx1_ASAP7_75t_R port map( A => n54, Y => n40);
   U59 : INVx1_ASAP7_75t_R port map( A => req(2), Y => n41);
   U60 : INVx1_ASAP7_75t_R port map( A => req(3), Y => n42);
   U61 : INVx1_ASAP7_75t_R port map( A => req(4), Y => n43);
   U62 : INVx1_ASAP7_75t_R port map( A => req(5), Y => n44);
   U63 : INVx1_ASAP7_75t_R port map( A => ack, Y => n45);
   U64 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n46);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT6_1 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (5 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (5 downto 0));

end rr_arbiter_no_delay_CNT6_1;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT6_1 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AO21x1_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI31xp33_ASAP7_75t_R
      port( A1, A2, A3, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OR3x1_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO32x1_ASAP7_75t_R
      port( A1, A2, A3, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_5_port, grant_4_port, grant_3_port, grant_2_port, grant_1_port,
      grant_0_port, pre_req_5_port, pre_req_4_port, pre_req_3_port, 
      pre_req_2_port, pre_req_1_port, pre_req_0_port, N2, N3, N4, N5, N6, 
      mask_pre_5_port, mask_pre_4_port, mask_pre_3_port, mask_pre_2_port, N20, 
      n1, n2_port, n3_port, n4_port, n5_port, n8, n9, n10, n11, n12, n13, n15, 
      n17, n19, n21, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
      n50, n51, n52, n53, n54, n55 : std_logic;

begin
   grant <= ( grant_5_port, grant_4_port, grant_3_port, grant_2_port, 
      grant_1_port, grant_0_port );
   
   U13 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(5), A3 => n4_port, 
                           B1 => n1, B2 => mask_pre_5_port, Y => grant_5_port);
   U14 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(4), A3 => n9, B1 => 
                           n21, B2 => mask_pre_4_port, Y => grant_4_port);
   U15 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(3), A3 => n5_port, 
                           B1 => n19, B2 => mask_pre_3_port, Y => grant_3_port)
                           ;
   U16 : AO32x1_ASAP7_75t_R port map( A1 => n55, A2 => req(2), A3 => n8, B1 => 
                           n17, B2 => mask_pre_2_port, Y => grant_2_port);
   U20 : OR3x1_ASAP7_75t_R port map( A => mask_pre_3_port, B => mask_pre_5_port
                           , C => mask_pre_4_port, Y => n54);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_4_port, A2 => ack, B1 => 
                           grant_4_port, B2 => n46, Y => n53);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_3_port, A2 => ack, B1 => 
                           grant_3_port, B2 => n46, Y => n52);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_2_port, A2 => ack, B1 => 
                           grant_2_port, B2 => n46, Y => n51);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_5_port, A2 => ack, B1 => 
                           grant_5_port, B2 => n46, Y => n50);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n46, Y => n49);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n46, Y => n48);
   pre_req_reg_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_4_port);
   pre_req_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n52, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_3_port);
   pre_req_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_2_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n49, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_1_port);
   pre_req_reg_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n50, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_5_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n48, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_0_port);
   U4 : TIELOx1_ASAP7_75t_R port map( L => n23);
   U5 : XOR2xp5_ASAP7_75t_R port map( A => n33, B => n15, Y => n1);
   U11 : AND2x2_ASAP7_75t_R port map( A => n41, B => n11, Y => n2_port);
   U12 : AND2x2_ASAP7_75t_R port map( A => n39, B => n10, Y => n3_port);
   U17 : XOR2xp5_ASAP7_75t_R port map( A => n45, B => n3_port, Y => n4_port);
   U18 : XOR2xp5_ASAP7_75t_R port map( A => n40, B => n2_port, Y => n5_port);
   U19 : XOR2xp5_ASAP7_75t_R port map( A => n41, B => n11, Y => n8);
   U21 : XOR2xp5_ASAP7_75t_R port map( A => n39, B => n10, Y => n9);
   U22 : AND2x2_ASAP7_75t_R port map( A => n40, B => n2_port, Y => n10);
   U23 : AND2x2_ASAP7_75t_R port map( A => n42, B => n43, Y => n11);
   U24 : AND2x2_ASAP7_75t_R port map( A => n36, B => n37, Y => n12);
   U25 : AND2x2_ASAP7_75t_R port map( A => n35, B => n12, Y => n13);
   U26 : AND2x2_ASAP7_75t_R port map( A => n34, B => n13, Y => n15);
   U27 : XOR2xp5_ASAP7_75t_R port map( A => n36, B => n37, Y => n17);
   U28 : XOR2xp5_ASAP7_75t_R port map( A => n35, B => n12, Y => n19);
   U29 : XOR2xp5_ASAP7_75t_R port map( A => n34, B => n13, Y => n21);
   U30 : NOR2xp33_ASAP7_75t_R port map( A => n44, B => n43, Y => grant_0_port);
   U31 : NOR3xp33_ASAP7_75t_R port map( A => n54, B => N20, C => 
                           mask_pre_2_port, Y => n55);
   U32 : INVx1_ASAP7_75t_R port map( A => rst, Y => n25);
   U33 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_5_port, B => N6, C => n45,
                           Y => mask_pre_5_port);
   U34 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_2_port, B => N3, C => n41,
                           Y => mask_pre_2_port);
   U35 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_1_port, B => N2, C => n47,
                           Y => N20);
   U36 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_4_port, B => N5, C => n39,
                           Y => mask_pre_4_port);
   U37 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_3_port, B => N4, C => n40,
                           Y => mask_pre_3_port);
   U38 : OAI31xp33_ASAP7_75t_R port map( A1 => n44, A2 => n38, A3 => n47, B => 
                           n37, Y => grant_1_port);
   U39 : XNOR2xp5_ASAP7_75t_R port map( A => n42, B => n43, Y => n38);
   U40 : NOR2xp33_ASAP7_75t_R port map( A => pre_req_1_port, B => 
                           pre_req_0_port, Y => n26);
   U41 : AO21x1_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => 
                           pre_req_1_port, B => n26, Y => N2);
   U42 : NOR2xp33_ASAP7_75t_R port map( A => n30, B => pre_req_2_port, Y => n27
                           );
   U43 : AO21x1_ASAP7_75t_R port map( A1 => n30, A2 => pre_req_2_port, B => n27
                           , Y => N3);
   U44 : NOR2xp33_ASAP7_75t_R port map( A => n31, B => pre_req_3_port, Y => n28
                           );
   U45 : AO21x1_ASAP7_75t_R port map( A1 => n31, A2 => pre_req_3_port, B => n28
                           , Y => N4);
   U46 : XNOR2xp5_ASAP7_75t_R port map( A => pre_req_4_port, B => n32, Y => N5)
                           ;
   U47 : NOR2xp33_ASAP7_75t_R port map( A => pre_req_4_port, B => n32, Y => n29
                           );
   U48 : XOR2xp5_ASAP7_75t_R port map( A => pre_req_5_port, B => n29, Y => N6);
   U49 : INVx1_ASAP7_75t_R port map( A => n26, Y => n30);
   U50 : INVx1_ASAP7_75t_R port map( A => n27, Y => n31);
   U51 : INVx1_ASAP7_75t_R port map( A => n28, Y => n32);
   U52 : INVx1_ASAP7_75t_R port map( A => mask_pre_5_port, Y => n33);
   U53 : INVx1_ASAP7_75t_R port map( A => mask_pre_4_port, Y => n34);
   U54 : INVx1_ASAP7_75t_R port map( A => mask_pre_3_port, Y => n35);
   U55 : INVx1_ASAP7_75t_R port map( A => mask_pre_2_port, Y => n36);
   U56 : INVx1_ASAP7_75t_R port map( A => N20, Y => n37);
   U57 : INVx1_ASAP7_75t_R port map( A => req(4), Y => n39);
   U58 : INVx1_ASAP7_75t_R port map( A => req(3), Y => n40);
   U59 : INVx1_ASAP7_75t_R port map( A => req(2), Y => n41);
   U60 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n42);
   U61 : INVx1_ASAP7_75t_R port map( A => req(0), Y => n43);
   U62 : INVx1_ASAP7_75t_R port map( A => n55, Y => n44);
   U63 : INVx1_ASAP7_75t_R port map( A => req(5), Y => n45);
   U64 : INVx1_ASAP7_75t_R port map( A => ack, Y => n46);
   U65 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n47);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity seq_packet_counter_1_12 is

   port( clk, rst, allocated : in std_logic;  packet_len : in std_logic_vector 
         (3 downto 0);  enr_vc : in std_logic;  flit_count : out 
         std_logic_vector (3 downto 0));

end seq_packet_counter_1_12;

architecture SYN_rtl of seq_packet_counter_1_12 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI311xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, C1 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13
      , n14, n15, n25, n26, n27, n28, n29, n30, n31, n32, n33 : std_logic;

begin
   flit_count <= ( flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port );
   
   U11 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(3), B => n30, Y => n31)
                           ;
   U12 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(2), B => n30, Y => n28)
                           ;
   U13 : OAI21xp5_ASAP7_75t_R port map( A1 => n30, A2 => n11, B => n27, Y => 
                           n29);
   U14 : NAND2xp5_ASAP7_75t_R port map( A => n26, B => n11, Y => n33);
   U15 : AOI21xp5_ASAP7_75t_R port map( A1 => n8, A2 => flit_count_0_port, B =>
                           n25, Y => n27);
   U26 : OAI311xp33_ASAP7_75t_R port map( A1 => n33, A2 => flit_count_3_port, 
                           A3 => flit_count_2_port, B1 => n32, C1 => n31, Y => 
                           n15);
   U27 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n8, B
                           => n29, C => flit_count_3_port, Y => n32);
   U28 : OAI221xp5_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n33, B1
                           => n7, B2 => n12, C => n28, Y => n14);
   U29 : OAI221xp5_ASAP7_75t_R port map( A1 => n10, A2 => n8, B1 => n11, B2 => 
                           n27, C => n33, Y => n13);
   flit_count_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_0_port);
   flit_count_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_1_port);
   flit_count_int_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_2_port);
   flit_count_int_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n5, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_3_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n2);
   U4 : AOI221xp5_ASAP7_75t_R port map( A1 => packet_len(0), A2 => n30, B1 => 
                           n25, B2 => flit_count_0_port, C => n26, Y => n1);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => enr_vc, Y => n30);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => enr_vc, B => allocated, Y => n25);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n3);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => n30, B => flit_count_0_port, C => 
                           n25, Y => n26);
   U9 : INVx1_ASAP7_75t_R port map( A => n13, Y => n4);
   U10 : INVx1_ASAP7_75t_R port map( A => n15, Y => n5);
   U16 : INVx1_ASAP7_75t_R port map( A => n14, Y => n6);
   U17 : INVx1_ASAP7_75t_R port map( A => n29, Y => n7);
   U18 : INVx1_ASAP7_75t_R port map( A => n30, Y => n8);
   U19 : INVx1_ASAP7_75t_R port map( A => allocated, Y => n9);
   U20 : INVx1_ASAP7_75t_R port map( A => packet_len(1), Y => n10);
   U21 : INVx1_ASAP7_75t_R port map( A => flit_count_1_port, Y => n11);
   U22 : INVx1_ASAP7_75t_R port map( A => flit_count_2_port, Y => n12);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity seq_packet_counter_1_11 is

   port( clk, rst, allocated : in std_logic;  packet_len : in std_logic_vector 
         (3 downto 0);  enr_vc : in std_logic;  flit_count : out 
         std_logic_vector (3 downto 0));

end seq_packet_counter_1_11;

architecture SYN_rtl of seq_packet_counter_1_11 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI311xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, C1 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13
      , n14, n15, n25, n26, n27, n28, n29, n30, n31, n32, n33 : std_logic;

begin
   flit_count <= ( flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port );
   
   U11 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(3), B => n30, Y => n31)
                           ;
   U12 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(2), B => n30, Y => n28)
                           ;
   U13 : OAI21xp5_ASAP7_75t_R port map( A1 => n30, A2 => n11, B => n27, Y => 
                           n29);
   U14 : NAND2xp5_ASAP7_75t_R port map( A => n26, B => n11, Y => n33);
   U15 : AOI21xp5_ASAP7_75t_R port map( A1 => n8, A2 => flit_count_0_port, B =>
                           n25, Y => n27);
   U26 : OAI311xp33_ASAP7_75t_R port map( A1 => n33, A2 => flit_count_3_port, 
                           A3 => flit_count_2_port, B1 => n32, C1 => n31, Y => 
                           n15);
   U27 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n8, B
                           => n29, C => flit_count_3_port, Y => n32);
   U28 : OAI221xp5_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n33, B1
                           => n7, B2 => n12, C => n28, Y => n14);
   U29 : OAI221xp5_ASAP7_75t_R port map( A1 => n10, A2 => n8, B1 => n11, B2 => 
                           n27, C => n33, Y => n13);
   flit_count_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_0_port);
   flit_count_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_1_port);
   flit_count_int_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_2_port);
   flit_count_int_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n5, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_3_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n2);
   U4 : AOI221xp5_ASAP7_75t_R port map( A1 => packet_len(0), A2 => n30, B1 => 
                           n25, B2 => flit_count_0_port, C => n26, Y => n1);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => enr_vc, Y => n30);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => enr_vc, B => allocated, Y => n25);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n3);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => n30, B => flit_count_0_port, C => 
                           n25, Y => n26);
   U9 : INVx1_ASAP7_75t_R port map( A => n13, Y => n4);
   U10 : INVx1_ASAP7_75t_R port map( A => n15, Y => n5);
   U16 : INVx1_ASAP7_75t_R port map( A => n14, Y => n6);
   U17 : INVx1_ASAP7_75t_R port map( A => n29, Y => n7);
   U18 : INVx1_ASAP7_75t_R port map( A => n30, Y => n8);
   U19 : INVx1_ASAP7_75t_R port map( A => allocated, Y => n9);
   U20 : INVx1_ASAP7_75t_R port map( A => packet_len(1), Y => n10);
   U21 : INVx1_ASAP7_75t_R port map( A => flit_count_1_port, Y => n11);
   U22 : INVx1_ASAP7_75t_R port map( A => flit_count_2_port, Y => n12);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity seq_packet_counter_1_10 is

   port( clk, rst, allocated : in std_logic;  packet_len : in std_logic_vector 
         (3 downto 0);  enr_vc : in std_logic;  flit_count : out 
         std_logic_vector (3 downto 0));

end seq_packet_counter_1_10;

architecture SYN_rtl of seq_packet_counter_1_10 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI311xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, C1 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13
      , n14, n15, n25, n26, n27, n28, n29, n30, n31, n32, n33 : std_logic;

begin
   flit_count <= ( flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port );
   
   U11 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(3), B => n30, Y => n31)
                           ;
   U12 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(2), B => n30, Y => n28)
                           ;
   U13 : OAI21xp5_ASAP7_75t_R port map( A1 => n30, A2 => n11, B => n27, Y => 
                           n29);
   U14 : NAND2xp5_ASAP7_75t_R port map( A => n26, B => n11, Y => n33);
   U15 : AOI21xp5_ASAP7_75t_R port map( A1 => n8, A2 => flit_count_0_port, B =>
                           n25, Y => n27);
   U26 : OAI311xp33_ASAP7_75t_R port map( A1 => n33, A2 => flit_count_3_port, 
                           A3 => flit_count_2_port, B1 => n32, C1 => n31, Y => 
                           n15);
   U27 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n8, B
                           => n29, C => flit_count_3_port, Y => n32);
   U28 : OAI221xp5_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n33, B1
                           => n7, B2 => n12, C => n28, Y => n14);
   U29 : OAI221xp5_ASAP7_75t_R port map( A1 => n10, A2 => n8, B1 => n11, B2 => 
                           n27, C => n33, Y => n13);
   flit_count_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_0_port);
   flit_count_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_1_port);
   flit_count_int_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_2_port);
   flit_count_int_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n5, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_3_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n2);
   U4 : AOI221xp5_ASAP7_75t_R port map( A1 => packet_len(0), A2 => n30, B1 => 
                           n25, B2 => flit_count_0_port, C => n26, Y => n1);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => enr_vc, Y => n30);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => enr_vc, B => allocated, Y => n25);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n3);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => n30, B => flit_count_0_port, C => 
                           n25, Y => n26);
   U9 : INVx1_ASAP7_75t_R port map( A => n13, Y => n4);
   U10 : INVx1_ASAP7_75t_R port map( A => n15, Y => n5);
   U16 : INVx1_ASAP7_75t_R port map( A => n14, Y => n6);
   U17 : INVx1_ASAP7_75t_R port map( A => n29, Y => n7);
   U18 : INVx1_ASAP7_75t_R port map( A => n30, Y => n8);
   U19 : INVx1_ASAP7_75t_R port map( A => allocated, Y => n9);
   U20 : INVx1_ASAP7_75t_R port map( A => packet_len(1), Y => n10);
   U21 : INVx1_ASAP7_75t_R port map( A => flit_count_1_port, Y => n11);
   U22 : INVx1_ASAP7_75t_R port map( A => flit_count_2_port, Y => n12);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity seq_packet_counter_1_9 is

   port( clk, rst, allocated : in std_logic;  packet_len : in std_logic_vector 
         (3 downto 0);  enr_vc : in std_logic;  flit_count : out 
         std_logic_vector (3 downto 0));

end seq_packet_counter_1_9;

architecture SYN_rtl of seq_packet_counter_1_9 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI311xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, C1 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13
      , n14, n15, n25, n26, n27, n28, n29, n30, n31, n32, n33 : std_logic;

begin
   flit_count <= ( flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port );
   
   U11 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(3), B => n30, Y => n31)
                           ;
   U12 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(2), B => n30, Y => n28)
                           ;
   U13 : OAI21xp5_ASAP7_75t_R port map( A1 => n30, A2 => n11, B => n27, Y => 
                           n29);
   U14 : NAND2xp5_ASAP7_75t_R port map( A => n26, B => n11, Y => n33);
   U15 : AOI21xp5_ASAP7_75t_R port map( A1 => n8, A2 => flit_count_0_port, B =>
                           n25, Y => n27);
   U26 : OAI311xp33_ASAP7_75t_R port map( A1 => n33, A2 => flit_count_3_port, 
                           A3 => flit_count_2_port, B1 => n32, C1 => n31, Y => 
                           n15);
   U27 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n8, B
                           => n29, C => flit_count_3_port, Y => n32);
   U28 : OAI221xp5_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n33, B1
                           => n7, B2 => n12, C => n28, Y => n14);
   U29 : OAI221xp5_ASAP7_75t_R port map( A1 => n10, A2 => n8, B1 => n11, B2 => 
                           n27, C => n33, Y => n13);
   flit_count_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_0_port);
   flit_count_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_1_port);
   flit_count_int_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_2_port);
   flit_count_int_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n5, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_3_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n2);
   U4 : AOI221xp5_ASAP7_75t_R port map( A1 => packet_len(0), A2 => n30, B1 => 
                           n25, B2 => flit_count_0_port, C => n26, Y => n1);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => enr_vc, Y => n30);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => enr_vc, B => allocated, Y => n25);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n3);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => n30, B => flit_count_0_port, C => 
                           n25, Y => n26);
   U9 : INVx1_ASAP7_75t_R port map( A => n13, Y => n4);
   U10 : INVx1_ASAP7_75t_R port map( A => n15, Y => n5);
   U16 : INVx1_ASAP7_75t_R port map( A => n14, Y => n6);
   U17 : INVx1_ASAP7_75t_R port map( A => n29, Y => n7);
   U18 : INVx1_ASAP7_75t_R port map( A => n30, Y => n8);
   U19 : INVx1_ASAP7_75t_R port map( A => allocated, Y => n9);
   U20 : INVx1_ASAP7_75t_R port map( A => packet_len(1), Y => n10);
   U21 : INVx1_ASAP7_75t_R port map( A => flit_count_1_port, Y => n11);
   U22 : INVx1_ASAP7_75t_R port map( A => flit_count_2_port, Y => n12);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity seq_packet_counter_1_8 is

   port( clk, rst, allocated : in std_logic;  packet_len : in std_logic_vector 
         (3 downto 0);  enr_vc : in std_logic;  flit_count : out 
         std_logic_vector (3 downto 0));

end seq_packet_counter_1_8;

architecture SYN_rtl of seq_packet_counter_1_8 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI311xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, C1 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13
      , n14, n15, n25, n26, n27, n28, n29, n30, n31, n32, n33 : std_logic;

begin
   flit_count <= ( flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port );
   
   U11 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(3), B => n30, Y => n31)
                           ;
   U12 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(2), B => n30, Y => n28)
                           ;
   U13 : OAI21xp5_ASAP7_75t_R port map( A1 => n30, A2 => n11, B => n27, Y => 
                           n29);
   U14 : NAND2xp5_ASAP7_75t_R port map( A => n26, B => n11, Y => n33);
   U15 : AOI21xp5_ASAP7_75t_R port map( A1 => n8, A2 => flit_count_0_port, B =>
                           n25, Y => n27);
   U26 : OAI311xp33_ASAP7_75t_R port map( A1 => n33, A2 => flit_count_3_port, 
                           A3 => flit_count_2_port, B1 => n32, C1 => n31, Y => 
                           n15);
   U27 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n8, B
                           => n29, C => flit_count_3_port, Y => n32);
   U28 : OAI221xp5_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n33, B1
                           => n7, B2 => n12, C => n28, Y => n14);
   U29 : OAI221xp5_ASAP7_75t_R port map( A1 => n10, A2 => n8, B1 => n11, B2 => 
                           n27, C => n33, Y => n13);
   flit_count_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_0_port);
   flit_count_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_1_port);
   flit_count_int_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_2_port);
   flit_count_int_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n5, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_3_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n2);
   U4 : AOI221xp5_ASAP7_75t_R port map( A1 => packet_len(0), A2 => n30, B1 => 
                           n25, B2 => flit_count_0_port, C => n26, Y => n1);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => enr_vc, Y => n30);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => enr_vc, B => allocated, Y => n25);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n3);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => n30, B => flit_count_0_port, C => 
                           n25, Y => n26);
   U9 : INVx1_ASAP7_75t_R port map( A => n13, Y => n4);
   U10 : INVx1_ASAP7_75t_R port map( A => n15, Y => n5);
   U16 : INVx1_ASAP7_75t_R port map( A => n14, Y => n6);
   U17 : INVx1_ASAP7_75t_R port map( A => n29, Y => n7);
   U18 : INVx1_ASAP7_75t_R port map( A => n30, Y => n8);
   U19 : INVx1_ASAP7_75t_R port map( A => allocated, Y => n9);
   U20 : INVx1_ASAP7_75t_R port map( A => packet_len(1), Y => n10);
   U21 : INVx1_ASAP7_75t_R port map( A => flit_count_1_port, Y => n11);
   U22 : INVx1_ASAP7_75t_R port map( A => flit_count_2_port, Y => n12);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity seq_packet_counter_1_7 is

   port( clk, rst, allocated : in std_logic;  packet_len : in std_logic_vector 
         (3 downto 0);  enr_vc : in std_logic;  flit_count : out 
         std_logic_vector (3 downto 0));

end seq_packet_counter_1_7;

architecture SYN_rtl of seq_packet_counter_1_7 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI311xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, C1 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13
      , n14, n15, n25, n26, n27, n28, n29, n30, n31, n32, n33 : std_logic;

begin
   flit_count <= ( flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port );
   
   U11 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(3), B => n30, Y => n31)
                           ;
   U12 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(2), B => n30, Y => n28)
                           ;
   U13 : OAI21xp5_ASAP7_75t_R port map( A1 => n30, A2 => n11, B => n27, Y => 
                           n29);
   U14 : NAND2xp5_ASAP7_75t_R port map( A => n26, B => n11, Y => n33);
   U15 : AOI21xp5_ASAP7_75t_R port map( A1 => n8, A2 => flit_count_0_port, B =>
                           n25, Y => n27);
   U26 : OAI311xp33_ASAP7_75t_R port map( A1 => n33, A2 => flit_count_3_port, 
                           A3 => flit_count_2_port, B1 => n32, C1 => n31, Y => 
                           n15);
   U27 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n8, B
                           => n29, C => flit_count_3_port, Y => n32);
   U28 : OAI221xp5_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n33, B1
                           => n7, B2 => n12, C => n28, Y => n14);
   U29 : OAI221xp5_ASAP7_75t_R port map( A1 => n10, A2 => n8, B1 => n11, B2 => 
                           n27, C => n33, Y => n13);
   flit_count_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_0_port);
   flit_count_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_1_port);
   flit_count_int_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_2_port);
   flit_count_int_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n5, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_3_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n2);
   U4 : AOI221xp5_ASAP7_75t_R port map( A1 => packet_len(0), A2 => n30, B1 => 
                           n25, B2 => flit_count_0_port, C => n26, Y => n1);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => enr_vc, Y => n30);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => enr_vc, B => allocated, Y => n25);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n3);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => n30, B => flit_count_0_port, C => 
                           n25, Y => n26);
   U9 : INVx1_ASAP7_75t_R port map( A => n13, Y => n4);
   U10 : INVx1_ASAP7_75t_R port map( A => n15, Y => n5);
   U16 : INVx1_ASAP7_75t_R port map( A => n14, Y => n6);
   U17 : INVx1_ASAP7_75t_R port map( A => n29, Y => n7);
   U18 : INVx1_ASAP7_75t_R port map( A => n30, Y => n8);
   U19 : INVx1_ASAP7_75t_R port map( A => allocated, Y => n9);
   U20 : INVx1_ASAP7_75t_R port map( A => packet_len(1), Y => n10);
   U21 : INVx1_ASAP7_75t_R port map( A => flit_count_1_port, Y => n11);
   U22 : INVx1_ASAP7_75t_R port map( A => flit_count_2_port, Y => n12);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity seq_packet_counter_1_6 is

   port( clk, rst, allocated : in std_logic;  packet_len : in std_logic_vector 
         (3 downto 0);  enr_vc : in std_logic;  flit_count : out 
         std_logic_vector (3 downto 0));

end seq_packet_counter_1_6;

architecture SYN_rtl of seq_packet_counter_1_6 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI311xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, C1 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13
      , n14, n15, n25, n26, n27, n28, n29, n30, n31, n32, n33 : std_logic;

begin
   flit_count <= ( flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port );
   
   U11 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(3), B => n30, Y => n31)
                           ;
   U12 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(2), B => n30, Y => n28)
                           ;
   U13 : OAI21xp5_ASAP7_75t_R port map( A1 => n30, A2 => n11, B => n27, Y => 
                           n29);
   U14 : NAND2xp5_ASAP7_75t_R port map( A => n26, B => n11, Y => n33);
   U15 : AOI21xp5_ASAP7_75t_R port map( A1 => n8, A2 => flit_count_0_port, B =>
                           n25, Y => n27);
   U26 : OAI311xp33_ASAP7_75t_R port map( A1 => n33, A2 => flit_count_3_port, 
                           A3 => flit_count_2_port, B1 => n32, C1 => n31, Y => 
                           n15);
   U27 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n8, B
                           => n29, C => flit_count_3_port, Y => n32);
   U28 : OAI221xp5_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n33, B1
                           => n7, B2 => n12, C => n28, Y => n14);
   U29 : OAI221xp5_ASAP7_75t_R port map( A1 => n10, A2 => n8, B1 => n11, B2 => 
                           n27, C => n33, Y => n13);
   flit_count_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_0_port);
   flit_count_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_1_port);
   flit_count_int_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_2_port);
   flit_count_int_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n5, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_3_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n2);
   U4 : AOI221xp5_ASAP7_75t_R port map( A1 => packet_len(0), A2 => n30, B1 => 
                           n25, B2 => flit_count_0_port, C => n26, Y => n1);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => enr_vc, Y => n30);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => enr_vc, B => allocated, Y => n25);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n3);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => n30, B => flit_count_0_port, C => 
                           n25, Y => n26);
   U9 : INVx1_ASAP7_75t_R port map( A => n13, Y => n4);
   U10 : INVx1_ASAP7_75t_R port map( A => n15, Y => n5);
   U16 : INVx1_ASAP7_75t_R port map( A => n14, Y => n6);
   U17 : INVx1_ASAP7_75t_R port map( A => n29, Y => n7);
   U18 : INVx1_ASAP7_75t_R port map( A => n30, Y => n8);
   U19 : INVx1_ASAP7_75t_R port map( A => allocated, Y => n9);
   U20 : INVx1_ASAP7_75t_R port map( A => packet_len(1), Y => n10);
   U21 : INVx1_ASAP7_75t_R port map( A => flit_count_1_port, Y => n11);
   U22 : INVx1_ASAP7_75t_R port map( A => flit_count_2_port, Y => n12);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity seq_packet_counter_1_5 is

   port( clk, rst, allocated : in std_logic;  packet_len : in std_logic_vector 
         (3 downto 0);  enr_vc : in std_logic;  flit_count : out 
         std_logic_vector (3 downto 0));

end seq_packet_counter_1_5;

architecture SYN_rtl of seq_packet_counter_1_5 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI311xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, C1 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13
      , n14, n15, n25, n26, n27, n28, n29, n30, n31, n32, n33 : std_logic;

begin
   flit_count <= ( flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port );
   
   U11 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(3), B => n30, Y => n31)
                           ;
   U12 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(2), B => n30, Y => n28)
                           ;
   U13 : OAI21xp5_ASAP7_75t_R port map( A1 => n30, A2 => n11, B => n27, Y => 
                           n29);
   U14 : NAND2xp5_ASAP7_75t_R port map( A => n26, B => n11, Y => n33);
   U15 : AOI21xp5_ASAP7_75t_R port map( A1 => n8, A2 => flit_count_0_port, B =>
                           n25, Y => n27);
   U26 : OAI311xp33_ASAP7_75t_R port map( A1 => n33, A2 => flit_count_3_port, 
                           A3 => flit_count_2_port, B1 => n32, C1 => n31, Y => 
                           n15);
   U27 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n8, B
                           => n29, C => flit_count_3_port, Y => n32);
   U28 : OAI221xp5_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n33, B1
                           => n7, B2 => n12, C => n28, Y => n14);
   U29 : OAI221xp5_ASAP7_75t_R port map( A1 => n10, A2 => n8, B1 => n11, B2 => 
                           n27, C => n33, Y => n13);
   flit_count_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_0_port);
   flit_count_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_1_port);
   flit_count_int_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_2_port);
   flit_count_int_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n5, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_3_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n2);
   U4 : AOI221xp5_ASAP7_75t_R port map( A1 => packet_len(0), A2 => n30, B1 => 
                           n25, B2 => flit_count_0_port, C => n26, Y => n1);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => enr_vc, Y => n30);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => enr_vc, B => allocated, Y => n25);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n3);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => n30, B => flit_count_0_port, C => 
                           n25, Y => n26);
   U9 : INVx1_ASAP7_75t_R port map( A => n13, Y => n4);
   U10 : INVx1_ASAP7_75t_R port map( A => n15, Y => n5);
   U16 : INVx1_ASAP7_75t_R port map( A => n14, Y => n6);
   U17 : INVx1_ASAP7_75t_R port map( A => n29, Y => n7);
   U18 : INVx1_ASAP7_75t_R port map( A => n30, Y => n8);
   U19 : INVx1_ASAP7_75t_R port map( A => allocated, Y => n9);
   U20 : INVx1_ASAP7_75t_R port map( A => packet_len(1), Y => n10);
   U21 : INVx1_ASAP7_75t_R port map( A => flit_count_1_port, Y => n11);
   U22 : INVx1_ASAP7_75t_R port map( A => flit_count_2_port, Y => n12);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity seq_packet_counter_1_4 is

   port( clk, rst, allocated : in std_logic;  packet_len : in std_logic_vector 
         (3 downto 0);  enr_vc : in std_logic;  flit_count : out 
         std_logic_vector (3 downto 0));

end seq_packet_counter_1_4;

architecture SYN_rtl of seq_packet_counter_1_4 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI311xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, C1 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13
      , n14, n15, n25, n26, n27, n28, n29, n30, n31, n32, n33 : std_logic;

begin
   flit_count <= ( flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port );
   
   U11 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(3), B => n30, Y => n31)
                           ;
   U12 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(2), B => n30, Y => n28)
                           ;
   U13 : OAI21xp5_ASAP7_75t_R port map( A1 => n30, A2 => n11, B => n27, Y => 
                           n29);
   U14 : NAND2xp5_ASAP7_75t_R port map( A => n26, B => n11, Y => n33);
   U15 : AOI21xp5_ASAP7_75t_R port map( A1 => n8, A2 => flit_count_0_port, B =>
                           n25, Y => n27);
   U26 : OAI311xp33_ASAP7_75t_R port map( A1 => n33, A2 => flit_count_3_port, 
                           A3 => flit_count_2_port, B1 => n32, C1 => n31, Y => 
                           n15);
   U27 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n8, B
                           => n29, C => flit_count_3_port, Y => n32);
   U28 : OAI221xp5_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n33, B1
                           => n7, B2 => n12, C => n28, Y => n14);
   U29 : OAI221xp5_ASAP7_75t_R port map( A1 => n10, A2 => n8, B1 => n11, B2 => 
                           n27, C => n33, Y => n13);
   flit_count_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_0_port);
   flit_count_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_1_port);
   flit_count_int_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_2_port);
   flit_count_int_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n5, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_3_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n2);
   U4 : AOI221xp5_ASAP7_75t_R port map( A1 => packet_len(0), A2 => n30, B1 => 
                           n25, B2 => flit_count_0_port, C => n26, Y => n1);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => enr_vc, Y => n30);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => enr_vc, B => allocated, Y => n25);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n3);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => n30, B => flit_count_0_port, C => 
                           n25, Y => n26);
   U9 : INVx1_ASAP7_75t_R port map( A => n13, Y => n4);
   U10 : INVx1_ASAP7_75t_R port map( A => n15, Y => n5);
   U16 : INVx1_ASAP7_75t_R port map( A => n14, Y => n6);
   U17 : INVx1_ASAP7_75t_R port map( A => n29, Y => n7);
   U18 : INVx1_ASAP7_75t_R port map( A => n30, Y => n8);
   U19 : INVx1_ASAP7_75t_R port map( A => allocated, Y => n9);
   U20 : INVx1_ASAP7_75t_R port map( A => packet_len(1), Y => n10);
   U21 : INVx1_ASAP7_75t_R port map( A => flit_count_1_port, Y => n11);
   U22 : INVx1_ASAP7_75t_R port map( A => flit_count_2_port, Y => n12);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity seq_packet_counter_1_3 is

   port( clk, rst, allocated : in std_logic;  packet_len : in std_logic_vector 
         (3 downto 0);  enr_vc : in std_logic;  flit_count : out 
         std_logic_vector (3 downto 0));

end seq_packet_counter_1_3;

architecture SYN_rtl of seq_packet_counter_1_3 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI311xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, C1 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13
      , n14, n15, n25, n26, n27, n28, n29, n30, n31, n32, n33 : std_logic;

begin
   flit_count <= ( flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port );
   
   U11 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(3), B => n30, Y => n31)
                           ;
   U12 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(2), B => n30, Y => n28)
                           ;
   U13 : OAI21xp5_ASAP7_75t_R port map( A1 => n30, A2 => n11, B => n27, Y => 
                           n29);
   U14 : NAND2xp5_ASAP7_75t_R port map( A => n26, B => n11, Y => n33);
   U15 : AOI21xp5_ASAP7_75t_R port map( A1 => n8, A2 => flit_count_0_port, B =>
                           n25, Y => n27);
   U26 : OAI311xp33_ASAP7_75t_R port map( A1 => n33, A2 => flit_count_3_port, 
                           A3 => flit_count_2_port, B1 => n32, C1 => n31, Y => 
                           n15);
   U27 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n8, B
                           => n29, C => flit_count_3_port, Y => n32);
   U28 : OAI221xp5_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n33, B1
                           => n7, B2 => n12, C => n28, Y => n14);
   U29 : OAI221xp5_ASAP7_75t_R port map( A1 => n10, A2 => n8, B1 => n11, B2 => 
                           n27, C => n33, Y => n13);
   flit_count_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_0_port);
   flit_count_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_1_port);
   flit_count_int_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_2_port);
   flit_count_int_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n5, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_3_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n2);
   U4 : AOI221xp5_ASAP7_75t_R port map( A1 => packet_len(0), A2 => n30, B1 => 
                           n25, B2 => flit_count_0_port, C => n26, Y => n1);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => enr_vc, Y => n30);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => enr_vc, B => allocated, Y => n25);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n3);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => n30, B => flit_count_0_port, C => 
                           n25, Y => n26);
   U9 : INVx1_ASAP7_75t_R port map( A => n13, Y => n4);
   U10 : INVx1_ASAP7_75t_R port map( A => n15, Y => n5);
   U16 : INVx1_ASAP7_75t_R port map( A => n14, Y => n6);
   U17 : INVx1_ASAP7_75t_R port map( A => n29, Y => n7);
   U18 : INVx1_ASAP7_75t_R port map( A => n30, Y => n8);
   U19 : INVx1_ASAP7_75t_R port map( A => allocated, Y => n9);
   U20 : INVx1_ASAP7_75t_R port map( A => packet_len(1), Y => n10);
   U21 : INVx1_ASAP7_75t_R port map( A => flit_count_1_port, Y => n11);
   U22 : INVx1_ASAP7_75t_R port map( A => flit_count_2_port, Y => n12);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity seq_packet_counter_1_2 is

   port( clk, rst, allocated : in std_logic;  packet_len : in std_logic_vector 
         (3 downto 0);  enr_vc : in std_logic;  flit_count : out 
         std_logic_vector (3 downto 0));

end seq_packet_counter_1_2;

architecture SYN_rtl of seq_packet_counter_1_2 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI311xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, C1 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13
      , n14, n15, n25, n26, n27, n28, n29, n30, n31, n32, n33 : std_logic;

begin
   flit_count <= ( flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port );
   
   U11 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(3), B => n30, Y => n31)
                           ;
   U12 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(2), B => n30, Y => n28)
                           ;
   U13 : OAI21xp5_ASAP7_75t_R port map( A1 => n30, A2 => n11, B => n27, Y => 
                           n29);
   U14 : NAND2xp5_ASAP7_75t_R port map( A => n26, B => n11, Y => n33);
   U15 : AOI21xp5_ASAP7_75t_R port map( A1 => n8, A2 => flit_count_0_port, B =>
                           n25, Y => n27);
   U26 : OAI311xp33_ASAP7_75t_R port map( A1 => n33, A2 => flit_count_3_port, 
                           A3 => flit_count_2_port, B1 => n32, C1 => n31, Y => 
                           n15);
   U27 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n8, B
                           => n29, C => flit_count_3_port, Y => n32);
   U28 : OAI221xp5_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n33, B1
                           => n7, B2 => n12, C => n28, Y => n14);
   U29 : OAI221xp5_ASAP7_75t_R port map( A1 => n10, A2 => n8, B1 => n11, B2 => 
                           n27, C => n33, Y => n13);
   flit_count_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_0_port);
   flit_count_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_1_port);
   flit_count_int_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_2_port);
   flit_count_int_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n5, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_3_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n2);
   U4 : AOI221xp5_ASAP7_75t_R port map( A1 => packet_len(0), A2 => n30, B1 => 
                           n25, B2 => flit_count_0_port, C => n26, Y => n1);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => enr_vc, Y => n30);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => enr_vc, B => allocated, Y => n25);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n3);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => n30, B => flit_count_0_port, C => 
                           n25, Y => n26);
   U9 : INVx1_ASAP7_75t_R port map( A => n13, Y => n4);
   U10 : INVx1_ASAP7_75t_R port map( A => n15, Y => n5);
   U16 : INVx1_ASAP7_75t_R port map( A => n14, Y => n6);
   U17 : INVx1_ASAP7_75t_R port map( A => n29, Y => n7);
   U18 : INVx1_ASAP7_75t_R port map( A => n30, Y => n8);
   U19 : INVx1_ASAP7_75t_R port map( A => allocated, Y => n9);
   U20 : INVx1_ASAP7_75t_R port map( A => packet_len(1), Y => n10);
   U21 : INVx1_ASAP7_75t_R port map( A => flit_count_1_port, Y => n11);
   U22 : INVx1_ASAP7_75t_R port map( A => flit_count_2_port, Y => n12);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity seq_packet_counter_1_1 is

   port( clk, rst, allocated : in std_logic;  packet_len : in std_logic_vector 
         (3 downto 0);  enr_vc : in std_logic;  flit_count : out 
         std_logic_vector (3 downto 0));

end seq_packet_counter_1_1;

architecture SYN_rtl of seq_packet_counter_1_1 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI311xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, C1 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13
      , n14, n15, n25, n26, n27, n28, n29, n30, n31, n32, n33 : std_logic;

begin
   flit_count <= ( flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port );
   
   U11 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(3), B => n30, Y => n31)
                           ;
   U12 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(2), B => n30, Y => n28)
                           ;
   U13 : OAI21xp5_ASAP7_75t_R port map( A1 => n30, A2 => n11, B => n27, Y => 
                           n29);
   U14 : NAND2xp5_ASAP7_75t_R port map( A => n26, B => n11, Y => n33);
   U15 : AOI21xp5_ASAP7_75t_R port map( A1 => n8, A2 => flit_count_0_port, B =>
                           n25, Y => n27);
   U26 : OAI311xp33_ASAP7_75t_R port map( A1 => n33, A2 => flit_count_3_port, 
                           A3 => flit_count_2_port, B1 => n32, C1 => n31, Y => 
                           n15);
   U27 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n8, B
                           => n29, C => flit_count_3_port, Y => n32);
   U28 : OAI221xp5_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n33, B1
                           => n7, B2 => n12, C => n28, Y => n14);
   U29 : OAI221xp5_ASAP7_75t_R port map( A1 => n10, A2 => n8, B1 => n11, B2 => 
                           n27, C => n33, Y => n13);
   flit_count_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_0_port);
   flit_count_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_1_port);
   flit_count_int_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_2_port);
   flit_count_int_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n5, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_3_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n2);
   U4 : AOI221xp5_ASAP7_75t_R port map( A1 => packet_len(0), A2 => n30, B1 => 
                           n25, B2 => flit_count_0_port, C => n26, Y => n1);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => enr_vc, Y => n30);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => enr_vc, B => allocated, Y => n25);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n3);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => n30, B => flit_count_0_port, C => 
                           n25, Y => n26);
   U9 : INVx1_ASAP7_75t_R port map( A => n13, Y => n4);
   U10 : INVx1_ASAP7_75t_R port map( A => n15, Y => n5);
   U16 : INVx1_ASAP7_75t_R port map( A => n14, Y => n6);
   U17 : INVx1_ASAP7_75t_R port map( A => n29, Y => n7);
   U18 : INVx1_ASAP7_75t_R port map( A => n30, Y => n8);
   U19 : INVx1_ASAP7_75t_R port map( A => allocated, Y => n9);
   U20 : INVx1_ASAP7_75t_R port map( A => packet_len(1), Y => n10);
   U21 : INVx1_ASAP7_75t_R port map( A => flit_count_1_port, Y => n11);
   U22 : INVx1_ASAP7_75t_R port map( A => flit_count_2_port, Y => n12);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_6 is

   port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;  
         routing : out std_logic_vector (6 downto 0));

end routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_6;

architecture SYN_rtl of routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_6 is

   component dxyu_routing_Xis1_Yis1_Zis1_6
      port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;
            routing : out std_logic_vector (6 downto 0));
   end component;

begin
   
   dxyu_routing_1 : dxyu_routing_Xis1_Yis1_Zis1_6 port map( address(5) => 
                           address(5), address(4) => address(4), address(3) => 
                           address(3), address(2) => address(2), address(1) => 
                           address(1), address(0) => address(0), enable => 
                           enable, routing(6) => routing(6), routing(5) => 
                           routing(5), routing(4) => routing(4), routing(3) => 
                           routing(3), routing(2) => routing(2), routing(1) => 
                           routing(1), routing(0) => routing(0));

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_5 is

   port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;  
         routing : out std_logic_vector (6 downto 0));

end routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_5;

architecture SYN_rtl of routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_5 is

   component dxyu_routing_Xis1_Yis1_Zis1_5
      port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;
            routing : out std_logic_vector (6 downto 0));
   end component;

begin
   
   dxyu_routing_1 : dxyu_routing_Xis1_Yis1_Zis1_5 port map( address(5) => 
                           address(5), address(4) => address(4), address(3) => 
                           address(3), address(2) => address(2), address(1) => 
                           address(1), address(0) => address(0), enable => 
                           enable, routing(6) => routing(6), routing(5) => 
                           routing(5), routing(4) => routing(4), routing(3) => 
                           routing(3), routing(2) => routing(2), routing(1) => 
                           routing(1), routing(0) => routing(0));

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_4 is

   port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;  
         routing : out std_logic_vector (6 downto 0));

end routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_4;

architecture SYN_rtl of routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_4 is

   component dxyu_routing_Xis1_Yis1_Zis1_4
      port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;
            routing : out std_logic_vector (6 downto 0));
   end component;

begin
   
   dxyu_routing_1 : dxyu_routing_Xis1_Yis1_Zis1_4 port map( address(5) => 
                           address(5), address(4) => address(4), address(3) => 
                           address(3), address(2) => address(2), address(1) => 
                           address(1), address(0) => address(0), enable => 
                           enable, routing(6) => routing(6), routing(5) => 
                           routing(5), routing(4) => routing(4), routing(3) => 
                           routing(3), routing(2) => routing(2), routing(1) => 
                           routing(1), routing(0) => routing(0));

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_3 is

   port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;  
         routing : out std_logic_vector (6 downto 0));

end routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_3;

architecture SYN_rtl of routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_3 is

   component dxyu_routing_Xis1_Yis1_Zis1_3
      port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;
            routing : out std_logic_vector (6 downto 0));
   end component;

begin
   
   dxyu_routing_1 : dxyu_routing_Xis1_Yis1_Zis1_3 port map( address(5) => 
                           address(5), address(4) => address(4), address(3) => 
                           address(3), address(2) => address(2), address(1) => 
                           address(1), address(0) => address(0), enable => 
                           enable, routing(6) => routing(6), routing(5) => 
                           routing(5), routing(4) => routing(4), routing(3) => 
                           routing(3), routing(2) => routing(2), routing(1) => 
                           routing(1), routing(0) => routing(0));

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_2 is

   port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;  
         routing : out std_logic_vector (6 downto 0));

end routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_2;

architecture SYN_rtl of routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_2 is

   component dxyu_routing_Xis1_Yis1_Zis1_2
      port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;
            routing : out std_logic_vector (6 downto 0));
   end component;

begin
   
   dxyu_routing_1 : dxyu_routing_Xis1_Yis1_Zis1_2 port map( address(5) => 
                           address(5), address(4) => address(4), address(3) => 
                           address(3), address(2) => address(2), address(1) => 
                           address(1), address(0) => address(0), enable => 
                           enable, routing(6) => routing(6), routing(5) => 
                           routing(5), routing(4) => routing(4), routing(3) => 
                           routing(3), routing(2) => routing(2), routing(1) => 
                           routing(1), routing(0) => routing(0));

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_1 is

   port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;  
         routing : out std_logic_vector (6 downto 0));

end routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_1;

architecture SYN_rtl of routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_1 is

   component dxyu_routing_Xis1_Yis1_Zis1_1
      port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;
            routing : out std_logic_vector (6 downto 0));
   end component;

begin
   
   dxyu_routing_1 : dxyu_routing_Xis1_Yis1_Zis1_1 port map( address(5) => 
                           address(5), address(4) => address(4), address(3) => 
                           address(3), address(2) => address(2), address(1) => 
                           address(1), address(0) => address(0), enable => 
                           enable, routing(6) => routing(6), routing(5) => 
                           routing(5), routing(4) => routing(4), routing(3) => 
                           routing(3), routing(2) => routing(2), routing(1) => 
                           routing(1), routing(0) => routing(0));

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity credit_count_single_vc_depth_out2_12 is

   port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
         std_logic);

end credit_count_single_vc_depth_out2_12;

architecture SYN_rtl of credit_count_single_vc_depth_out2_12 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_val_1_port, count_val_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n13 : std_logic;

begin
   
   U10 : NAND2xp5_ASAP7_75t_R port map( A => vc_write_tx, B => n7, Y => n8);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => incr_rx, B => count_val_0_port, Y 
                           => n10);
   U15 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n5, A2 => n10, B => n9, C => 
                           n6, Y => n11);
   U16 : XNOR2xp5_ASAP7_75t_R port map( A => n10, B => n5, Y => n13);
   U17 : NAND3xp33_ASAP7_75t_R port map( A => n10, B => n6, C => n7, Y => 
                           credit_avail);
   U18 : XNOR2xp5_ASAP7_75t_R port map( A => count_val_0_port, B => incr_rx, Y 
                           => n7);
   count_val_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK => 
                           clk, RESET => n3, SET => n4, QN => count_val_1_port)
                           ;
   count_val_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2, CLK => 
                           clk, RESET => n4, SET => n3, QN => count_val_0_port)
                           ;
   U3 : TIELOx1_ASAP7_75t_R port map( L => n3);
   U4 : OA21x2_ASAP7_75t_R port map( A1 => n6, A2 => n13, B => n11, Y => n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => vc_write_tx, A2 => n7, B => n8, Y =>
                           n2);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx, B => n10, Y => n9);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n4);
   U8 : INVx1_ASAP7_75t_R port map( A => n8, Y => n5);
   U9 : INVx1_ASAP7_75t_R port map( A => count_val_1_port, Y => n6);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity credit_count_single_vc_depth_out2_11 is

   port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
         std_logic);

end credit_count_single_vc_depth_out2_11;

architecture SYN_rtl of credit_count_single_vc_depth_out2_11 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_val_1_port, count_val_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n13 : std_logic;

begin
   
   U10 : NAND2xp5_ASAP7_75t_R port map( A => vc_write_tx, B => n7, Y => n8);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => incr_rx, B => count_val_0_port, Y 
                           => n10);
   U15 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n5, A2 => n10, B => n9, C => 
                           n6, Y => n11);
   U16 : XNOR2xp5_ASAP7_75t_R port map( A => n10, B => n5, Y => n13);
   U17 : NAND3xp33_ASAP7_75t_R port map( A => n10, B => n6, C => n7, Y => 
                           credit_avail);
   U18 : XNOR2xp5_ASAP7_75t_R port map( A => count_val_0_port, B => incr_rx, Y 
                           => n7);
   count_val_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK => 
                           clk, RESET => n3, SET => n4, QN => count_val_1_port)
                           ;
   count_val_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2, CLK => 
                           clk, RESET => n4, SET => n3, QN => count_val_0_port)
                           ;
   U3 : TIELOx1_ASAP7_75t_R port map( L => n3);
   U4 : OA21x2_ASAP7_75t_R port map( A1 => n6, A2 => n13, B => n11, Y => n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => vc_write_tx, A2 => n7, B => n8, Y =>
                           n2);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx, B => n10, Y => n9);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n4);
   U8 : INVx1_ASAP7_75t_R port map( A => n8, Y => n5);
   U9 : INVx1_ASAP7_75t_R port map( A => count_val_1_port, Y => n6);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity credit_count_single_vc_depth_out2_10 is

   port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
         std_logic);

end credit_count_single_vc_depth_out2_10;

architecture SYN_rtl of credit_count_single_vc_depth_out2_10 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_val_1_port, count_val_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n13 : std_logic;

begin
   
   U10 : NAND2xp5_ASAP7_75t_R port map( A => vc_write_tx, B => n7, Y => n8);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => incr_rx, B => count_val_0_port, Y 
                           => n10);
   U15 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n5, A2 => n10, B => n9, C => 
                           n6, Y => n11);
   U16 : XNOR2xp5_ASAP7_75t_R port map( A => n10, B => n5, Y => n13);
   U17 : NAND3xp33_ASAP7_75t_R port map( A => n10, B => n6, C => n7, Y => 
                           credit_avail);
   U18 : XNOR2xp5_ASAP7_75t_R port map( A => count_val_0_port, B => incr_rx, Y 
                           => n7);
   count_val_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK => 
                           clk, RESET => n3, SET => n4, QN => count_val_1_port)
                           ;
   count_val_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2, CLK => 
                           clk, RESET => n4, SET => n3, QN => count_val_0_port)
                           ;
   U3 : TIELOx1_ASAP7_75t_R port map( L => n3);
   U4 : OA21x2_ASAP7_75t_R port map( A1 => n6, A2 => n13, B => n11, Y => n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => vc_write_tx, A2 => n7, B => n8, Y =>
                           n2);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx, B => n10, Y => n9);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n4);
   U8 : INVx1_ASAP7_75t_R port map( A => n8, Y => n5);
   U9 : INVx1_ASAP7_75t_R port map( A => count_val_1_port, Y => n6);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity credit_count_single_vc_depth_out2_9 is

   port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
         std_logic);

end credit_count_single_vc_depth_out2_9;

architecture SYN_rtl of credit_count_single_vc_depth_out2_9 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_val_1_port, count_val_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n13 : std_logic;

begin
   
   U10 : NAND2xp5_ASAP7_75t_R port map( A => vc_write_tx, B => n7, Y => n8);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => incr_rx, B => count_val_0_port, Y 
                           => n10);
   U15 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n5, A2 => n10, B => n9, C => 
                           n6, Y => n11);
   U16 : XNOR2xp5_ASAP7_75t_R port map( A => n10, B => n5, Y => n13);
   U17 : NAND3xp33_ASAP7_75t_R port map( A => n10, B => n6, C => n7, Y => 
                           credit_avail);
   U18 : XNOR2xp5_ASAP7_75t_R port map( A => count_val_0_port, B => incr_rx, Y 
                           => n7);
   count_val_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK => 
                           clk, RESET => n3, SET => n4, QN => count_val_1_port)
                           ;
   count_val_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2, CLK => 
                           clk, RESET => n4, SET => n3, QN => count_val_0_port)
                           ;
   U3 : TIELOx1_ASAP7_75t_R port map( L => n3);
   U4 : OA21x2_ASAP7_75t_R port map( A1 => n6, A2 => n13, B => n11, Y => n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => vc_write_tx, A2 => n7, B => n8, Y =>
                           n2);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx, B => n10, Y => n9);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n4);
   U8 : INVx1_ASAP7_75t_R port map( A => n8, Y => n5);
   U9 : INVx1_ASAP7_75t_R port map( A => count_val_1_port, Y => n6);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity credit_count_single_vc_depth_out2_8 is

   port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
         std_logic);

end credit_count_single_vc_depth_out2_8;

architecture SYN_rtl of credit_count_single_vc_depth_out2_8 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_val_1_port, count_val_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n13 : std_logic;

begin
   
   U10 : NAND2xp5_ASAP7_75t_R port map( A => vc_write_tx, B => n7, Y => n8);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => incr_rx, B => count_val_0_port, Y 
                           => n10);
   U15 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n5, A2 => n10, B => n9, C => 
                           n6, Y => n11);
   U16 : XNOR2xp5_ASAP7_75t_R port map( A => n10, B => n5, Y => n13);
   U17 : NAND3xp33_ASAP7_75t_R port map( A => n10, B => n6, C => n7, Y => 
                           credit_avail);
   U18 : XNOR2xp5_ASAP7_75t_R port map( A => count_val_0_port, B => incr_rx, Y 
                           => n7);
   count_val_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK => 
                           clk, RESET => n3, SET => n4, QN => count_val_1_port)
                           ;
   count_val_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2, CLK => 
                           clk, RESET => n4, SET => n3, QN => count_val_0_port)
                           ;
   U3 : TIELOx1_ASAP7_75t_R port map( L => n3);
   U4 : OA21x2_ASAP7_75t_R port map( A1 => n6, A2 => n13, B => n11, Y => n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => vc_write_tx, A2 => n7, B => n8, Y =>
                           n2);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx, B => n10, Y => n9);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n4);
   U8 : INVx1_ASAP7_75t_R port map( A => n8, Y => n5);
   U9 : INVx1_ASAP7_75t_R port map( A => count_val_1_port, Y => n6);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity credit_count_single_vc_depth_out2_7 is

   port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
         std_logic);

end credit_count_single_vc_depth_out2_7;

architecture SYN_rtl of credit_count_single_vc_depth_out2_7 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_val_1_port, count_val_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n13 : std_logic;

begin
   
   U10 : NAND2xp5_ASAP7_75t_R port map( A => vc_write_tx, B => n7, Y => n8);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => incr_rx, B => count_val_0_port, Y 
                           => n10);
   U15 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n5, A2 => n10, B => n9, C => 
                           n6, Y => n11);
   U16 : XNOR2xp5_ASAP7_75t_R port map( A => n10, B => n5, Y => n13);
   U17 : NAND3xp33_ASAP7_75t_R port map( A => n10, B => n6, C => n7, Y => 
                           credit_avail);
   U18 : XNOR2xp5_ASAP7_75t_R port map( A => count_val_0_port, B => incr_rx, Y 
                           => n7);
   count_val_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK => 
                           clk, RESET => n3, SET => n4, QN => count_val_1_port)
                           ;
   count_val_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2, CLK => 
                           clk, RESET => n4, SET => n3, QN => count_val_0_port)
                           ;
   U3 : TIELOx1_ASAP7_75t_R port map( L => n3);
   U4 : OA21x2_ASAP7_75t_R port map( A1 => n6, A2 => n13, B => n11, Y => n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => vc_write_tx, A2 => n7, B => n8, Y =>
                           n2);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx, B => n10, Y => n9);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n4);
   U8 : INVx1_ASAP7_75t_R port map( A => n8, Y => n5);
   U9 : INVx1_ASAP7_75t_R port map( A => count_val_1_port, Y => n6);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity credit_count_single_vc_depth_out2_6 is

   port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
         std_logic);

end credit_count_single_vc_depth_out2_6;

architecture SYN_rtl of credit_count_single_vc_depth_out2_6 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_val_1_port, count_val_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n13 : std_logic;

begin
   
   U10 : NAND2xp5_ASAP7_75t_R port map( A => vc_write_tx, B => n7, Y => n8);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => incr_rx, B => count_val_0_port, Y 
                           => n10);
   U15 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n5, A2 => n10, B => n9, C => 
                           n6, Y => n11);
   U16 : XNOR2xp5_ASAP7_75t_R port map( A => n10, B => n5, Y => n13);
   U17 : NAND3xp33_ASAP7_75t_R port map( A => n10, B => n6, C => n7, Y => 
                           credit_avail);
   U18 : XNOR2xp5_ASAP7_75t_R port map( A => count_val_0_port, B => incr_rx, Y 
                           => n7);
   count_val_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK => 
                           clk, RESET => n3, SET => n4, QN => count_val_1_port)
                           ;
   count_val_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2, CLK => 
                           clk, RESET => n4, SET => n3, QN => count_val_0_port)
                           ;
   U3 : TIELOx1_ASAP7_75t_R port map( L => n3);
   U4 : OA21x2_ASAP7_75t_R port map( A1 => n6, A2 => n13, B => n11, Y => n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => vc_write_tx, A2 => n7, B => n8, Y =>
                           n2);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx, B => n10, Y => n9);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n4);
   U8 : INVx1_ASAP7_75t_R port map( A => n8, Y => n5);
   U9 : INVx1_ASAP7_75t_R port map( A => count_val_1_port, Y => n6);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity credit_count_single_vc_depth_out2_5 is

   port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
         std_logic);

end credit_count_single_vc_depth_out2_5;

architecture SYN_rtl of credit_count_single_vc_depth_out2_5 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_val_1_port, count_val_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n13 : std_logic;

begin
   
   U10 : NAND2xp5_ASAP7_75t_R port map( A => vc_write_tx, B => n7, Y => n8);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => incr_rx, B => count_val_0_port, Y 
                           => n10);
   U15 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n5, A2 => n10, B => n9, C => 
                           n6, Y => n11);
   U16 : XNOR2xp5_ASAP7_75t_R port map( A => n10, B => n5, Y => n13);
   U17 : NAND3xp33_ASAP7_75t_R port map( A => n10, B => n6, C => n7, Y => 
                           credit_avail);
   U18 : XNOR2xp5_ASAP7_75t_R port map( A => count_val_0_port, B => incr_rx, Y 
                           => n7);
   count_val_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK => 
                           clk, RESET => n3, SET => n4, QN => count_val_1_port)
                           ;
   count_val_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2, CLK => 
                           clk, RESET => n4, SET => n3, QN => count_val_0_port)
                           ;
   U3 : TIELOx1_ASAP7_75t_R port map( L => n3);
   U4 : OA21x2_ASAP7_75t_R port map( A1 => n6, A2 => n13, B => n11, Y => n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => vc_write_tx, A2 => n7, B => n8, Y =>
                           n2);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx, B => n10, Y => n9);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n4);
   U8 : INVx1_ASAP7_75t_R port map( A => n8, Y => n5);
   U9 : INVx1_ASAP7_75t_R port map( A => count_val_1_port, Y => n6);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity credit_count_single_vc_depth_out2_4 is

   port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
         std_logic);

end credit_count_single_vc_depth_out2_4;

architecture SYN_rtl of credit_count_single_vc_depth_out2_4 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_val_1_port, count_val_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n13 : std_logic;

begin
   
   U10 : NAND2xp5_ASAP7_75t_R port map( A => vc_write_tx, B => n7, Y => n8);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => incr_rx, B => count_val_0_port, Y 
                           => n10);
   U15 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n5, A2 => n10, B => n9, C => 
                           n6, Y => n11);
   U16 : XNOR2xp5_ASAP7_75t_R port map( A => n10, B => n5, Y => n13);
   U17 : NAND3xp33_ASAP7_75t_R port map( A => n10, B => n6, C => n7, Y => 
                           credit_avail);
   U18 : XNOR2xp5_ASAP7_75t_R port map( A => count_val_0_port, B => incr_rx, Y 
                           => n7);
   count_val_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK => 
                           clk, RESET => n3, SET => n4, QN => count_val_1_port)
                           ;
   count_val_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2, CLK => 
                           clk, RESET => n4, SET => n3, QN => count_val_0_port)
                           ;
   U3 : TIELOx1_ASAP7_75t_R port map( L => n3);
   U4 : OA21x2_ASAP7_75t_R port map( A1 => n6, A2 => n13, B => n11, Y => n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => vc_write_tx, A2 => n7, B => n8, Y =>
                           n2);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx, B => n10, Y => n9);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n4);
   U8 : INVx1_ASAP7_75t_R port map( A => n8, Y => n5);
   U9 : INVx1_ASAP7_75t_R port map( A => count_val_1_port, Y => n6);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity credit_count_single_vc_depth_out2_3 is

   port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
         std_logic);

end credit_count_single_vc_depth_out2_3;

architecture SYN_rtl of credit_count_single_vc_depth_out2_3 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_val_1_port, count_val_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n13 : std_logic;

begin
   
   U10 : NAND2xp5_ASAP7_75t_R port map( A => vc_write_tx, B => n7, Y => n8);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => incr_rx, B => count_val_0_port, Y 
                           => n10);
   U15 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n5, A2 => n10, B => n9, C => 
                           n6, Y => n11);
   U16 : XNOR2xp5_ASAP7_75t_R port map( A => n10, B => n5, Y => n13);
   U17 : NAND3xp33_ASAP7_75t_R port map( A => n10, B => n6, C => n7, Y => 
                           credit_avail);
   U18 : XNOR2xp5_ASAP7_75t_R port map( A => count_val_0_port, B => incr_rx, Y 
                           => n7);
   count_val_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK => 
                           clk, RESET => n3, SET => n4, QN => count_val_1_port)
                           ;
   count_val_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2, CLK => 
                           clk, RESET => n4, SET => n3, QN => count_val_0_port)
                           ;
   U3 : TIELOx1_ASAP7_75t_R port map( L => n3);
   U4 : OA21x2_ASAP7_75t_R port map( A1 => n6, A2 => n13, B => n11, Y => n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => vc_write_tx, A2 => n7, B => n8, Y =>
                           n2);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx, B => n10, Y => n9);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n4);
   U8 : INVx1_ASAP7_75t_R port map( A => n8, Y => n5);
   U9 : INVx1_ASAP7_75t_R port map( A => count_val_1_port, Y => n6);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity credit_count_single_vc_depth_out2_2 is

   port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
         std_logic);

end credit_count_single_vc_depth_out2_2;

architecture SYN_rtl of credit_count_single_vc_depth_out2_2 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_val_1_port, count_val_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n13 : std_logic;

begin
   
   U10 : NAND2xp5_ASAP7_75t_R port map( A => vc_write_tx, B => n7, Y => n8);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => incr_rx, B => count_val_0_port, Y 
                           => n10);
   U15 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n5, A2 => n10, B => n9, C => 
                           n6, Y => n11);
   U16 : XNOR2xp5_ASAP7_75t_R port map( A => n10, B => n5, Y => n13);
   U17 : NAND3xp33_ASAP7_75t_R port map( A => n10, B => n6, C => n7, Y => 
                           credit_avail);
   U18 : XNOR2xp5_ASAP7_75t_R port map( A => count_val_0_port, B => incr_rx, Y 
                           => n7);
   count_val_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK => 
                           clk, RESET => n3, SET => n4, QN => count_val_1_port)
                           ;
   count_val_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2, CLK => 
                           clk, RESET => n4, SET => n3, QN => count_val_0_port)
                           ;
   U3 : TIELOx1_ASAP7_75t_R port map( L => n3);
   U4 : OA21x2_ASAP7_75t_R port map( A1 => n6, A2 => n13, B => n11, Y => n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => vc_write_tx, A2 => n7, B => n8, Y =>
                           n2);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx, B => n10, Y => n9);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n4);
   U8 : INVx1_ASAP7_75t_R port map( A => n8, Y => n5);
   U9 : INVx1_ASAP7_75t_R port map( A => count_val_1_port, Y => n6);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity credit_count_single_vc_depth_out2_1 is

   port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
         std_logic);

end credit_count_single_vc_depth_out2_1;

architecture SYN_rtl of credit_count_single_vc_depth_out2_1 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_val_1_port, count_val_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n13 : std_logic;

begin
   
   U10 : NAND2xp5_ASAP7_75t_R port map( A => vc_write_tx, B => n7, Y => n8);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => incr_rx, B => count_val_0_port, Y 
                           => n10);
   U15 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n5, A2 => n10, B => n9, C => 
                           n6, Y => n11);
   U16 : XNOR2xp5_ASAP7_75t_R port map( A => n10, B => n5, Y => n13);
   U17 : NAND3xp33_ASAP7_75t_R port map( A => n10, B => n6, C => n7, Y => 
                           credit_avail);
   U18 : XNOR2xp5_ASAP7_75t_R port map( A => count_val_0_port, B => incr_rx, Y 
                           => n7);
   count_val_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK => 
                           clk, RESET => n3, SET => n4, QN => count_val_1_port)
                           ;
   count_val_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2, CLK => 
                           clk, RESET => n4, SET => n3, QN => count_val_0_port)
                           ;
   U3 : TIELOx1_ASAP7_75t_R port map( L => n3);
   U4 : OA21x2_ASAP7_75t_R port map( A1 => n6, A2 => n13, B => n11, Y => n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => vc_write_tx, A2 => n7, B => n8, Y =>
                           n2);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx, B => n10, Y => n9);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n4);
   U8 : INVx1_ASAP7_75t_R port map( A => n8, Y => n5);
   U9 : INVx1_ASAP7_75t_R port map( A => count_val_1_port, Y => n6);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_17 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_17;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_17 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n5, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n3, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n3, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n4, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => ack, Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_16 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_16;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_16 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n5, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n3, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n3, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n4, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => ack, Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_15 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_15;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_15 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n5, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n3, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n3, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n4, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => ack, Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_14 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_14;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_14 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n5, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n3, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n3, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n4, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => ack, Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_13 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_13;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_13 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n5, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n3, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n3, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n4, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => ack, Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_12 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_12;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_12 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n4, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n5, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n5, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n3, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => ack, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_11 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_11;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_11 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n4, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n5, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n5, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n3, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => ack, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_10 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_10;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_10 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n4, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n5, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n5, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n3, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => ack, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_9 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_9;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_9 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n4, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n5, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n5, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n3, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => ack, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_8 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_8;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_8 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n4, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n5, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n5, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n3, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => ack, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_7 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_7;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_7 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n4, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n5, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n5, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n3, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => ack, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_6 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_6;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_6 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n5, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n3, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n3, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n4, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => ack, Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_5 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_5;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_5 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n5, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n3, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n3, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n4, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => ack, Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_4 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_4;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_4 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n5, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n3, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n3, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n4, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => ack, Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_3 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_3;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_3 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n5, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n3, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n3, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n4, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => ack, Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_2 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_2;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_2 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n5, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n3, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n3, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n4, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => ack, Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_1 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_1;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_1 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n1, n2, 
      n3, n4, n5, n6, n8, n9 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n9, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n5, C => 
                           pre_req_0_port, Y => n9);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n3, Y => n8);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n3, Y => n6);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n4, B => n9, Y => 
                           grant_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_0_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => ack, Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity vc_output_allocator_port_num7_vc_num_out2_5 is

   port( clk, rst : in std_logic;  rq_vc_out : in std_logic_vector (5 downto 0)
         ;  granted_vc, packet_end : in std_logic_vector (11 downto 0);  
         crossbar_ctrl_vec : out std_logic_vector (5 downto 0);  vc_sel_enc, 
         output_vc_in_use : out std_logic_vector (1 downto 0);  ack_rq_vc_out :
         out std_logic_vector (5 downto 0));

end vc_output_allocator_port_num7_vc_num_out2_5;

architecture SYN_rtl of vc_output_allocator_port_num7_vc_num_out2_5 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component rr_arbiter_no_delay_CNT6_5
      port( clk, rst : in std_logic;  req : in std_logic_vector (5 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (5 downto 0));
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI211xp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OA211x2_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1O1Ixp25_ASAP7_75t_R
      port( A1, A2, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal crossbar_ctrl_vec_5_port, crossbar_ctrl_vec_4_port, n124, 
      crossbar_ctrl_vec_2_port, crossbar_ctrl_vec_1_port, n125, 
      vc_sel_enc_1_0_port, vc_sel_enc_0_0_port, output_vc_in_use_1_port, 
      output_vc_in_use_0_port, vc_available, grant_5_port, grant_4_port, 
      grant_3_port, grant_2_port, grant_1_port, grant_0_port, n1, n2, n3, n4, 
      n5, crossbar_ctrl_vec_3_port, crossbar_ctrl_vec_0_port, n8, n9, n10, n11,
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123 : std_logic;

begin
   crossbar_ctrl_vec <= ( crossbar_ctrl_vec_5_port, crossbar_ctrl_vec_4_port, 
      crossbar_ctrl_vec_3_port, crossbar_ctrl_vec_2_port, 
      crossbar_ctrl_vec_1_port, crossbar_ctrl_vec_0_port );
   vc_sel_enc <= ( vc_sel_enc_1_0_port, vc_sel_enc_0_0_port );
   output_vc_in_use <= ( output_vc_in_use_1_port, output_vc_in_use_0_port );
   
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => n123, A2 => n13, B1 => n122, B2 
                           => n27, Y => n38);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => n121, A2 => n13, B1 => n122, B2 
                           => n28, Y => n37);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => n120, A2 => n13, B1 => n122, B2 
                           => n29, Y => n36);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => n123, A2 => n16, B1 => n119, B2 
                           => n23, Y => n35);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => n121, A2 => n16, B1 => n119, B2 
                           => n24, Y => n34);
   U28 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n116, A2 => n115, B => n25, C 
                           => n114, Y => n117);
   U30 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n30, B => n110, C => vc_sel_enc_0_0_port, Y => n111)
                           ;
   U31 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(2), B => 
                           crossbar_ctrl_vec_0_port, Y => n110);
   U33 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n22, B => n109, C => n24, Y => n115);
   U34 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(10), B => 
                           crossbar_ctrl_vec_0_port, Y => n109);
   U35 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n20, B => n108, C => n23, Y => n116);
   U36 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(6), B => 
                           crossbar_ctrl_vec_0_port, Y => n108);
   U37 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n107, A2 => n106, B => 
                           vc_sel_enc_0_0_port, C => n26, Y => n118);
   U38 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n32, B => n105, C => n24, Y => n106);
   U39 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(11), B => 
                           crossbar_ctrl_vec_0_port, Y => n105);
   U40 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n21, B => n104, C => n23, Y => n107);
   U41 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(7), B => 
                           crossbar_ctrl_vec_0_port, Y => n104);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => n120, A2 => n16, B1 => n119, B2 
                           => n25, Y => n33);
   U52 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_3_port, A2 =>
                           n31, B => n84, C => n29, Y => n85);
   U53 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(3), B => 
                           crossbar_ctrl_vec_3_port, Y => n84);
   U54 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_3_port, A2 =>
                           n30, B => n83, C => vc_sel_enc_1_0_port, Y => n86);
   U55 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(2), B => 
                           crossbar_ctrl_vec_3_port, Y => n83);
   U58 : NAND2xp5_ASAP7_75t_R port map( A => output_vc_in_use_1_port, B => 
                           output_vc_in_use_0_port, Y => vc_available);
   U81 : A2O1A1O1Ixp25_ASAP7_75t_R port map( A1 => packet_end(3), A2 => 
                           crossbar_ctrl_vec_0_port, B => n112, C => 
                           vc_sel_enc_0_0_port, D => n111, Y => n113);
   U82 : OA211x2_ASAP7_75t_R port map( A1 => n19, A2 => n102, B => n101, C => 
                           n100, Y => n120);
   U83 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(9), A2 => n99, B =>
                           n98, C => n18, Y => n100);
   U84 : AND2x2_ASAP7_75t_R port map( A => granted_vc(11), B => n17, Y => n98);
   U85 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(5), A2 => n99, B =>
                           n97, C => n19, Y => n101);
   U86 : AND2x2_ASAP7_75t_R port map( A => granted_vc(7), B => n17, Y => n97);
   U87 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(1), A2 => n99, B =>
                           n96, C => n121, Y => n102);
   U88 : AND2x2_ASAP7_75t_R port map( A => granted_vc(3), B => n17, Y => n96);
   U89 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n93, A2 => n92, B => n29, C =>
                           output_vc_in_use_1_port, Y => n94);
   U90 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(7), A2 => 
                           crossbar_ctrl_vec_3_port, B => n91, C => 
                           crossbar_ctrl_vec_4_port, Y => n92);
   U91 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(11), A2 => 
                           crossbar_ctrl_vec_3_port, B => n90, C => 
                           crossbar_ctrl_vec_5_port, Y => n93);
   U92 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n89, A2 => n88, B => 
                           vc_sel_enc_1_0_port, C => n87, Y => n95);
   U93 : OAI211xp5_ASAP7_75t_R port map( A1 => n86, A2 => n85, B => n27, C => 
                           n28, Y => n87);
   U94 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(6), A2 => 
                           crossbar_ctrl_vec_3_port, B => n82, C => 
                           crossbar_ctrl_vec_4_port, Y => n88);
   U95 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(10), A2 => 
                           crossbar_ctrl_vec_3_port, B => n39, C => 
                           crossbar_ctrl_vec_5_port, Y => n89);
   U96 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_5_port, Y 
                           => ack_rq_vc_out(5));
   U97 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_4_port, Y 
                           => ack_rq_vc_out(4));
   U98 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_3_port, Y 
                           => ack_rq_vc_out(3));
   U99 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_2_port, Y 
                           => ack_rq_vc_out(2));
   U100 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_1_port, Y 
                           => ack_rq_vc_out(1));
   U101 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_0_port, Y 
                           => ack_rq_vc_out(0));
   rr_arbiter : rr_arbiter_no_delay_CNT6_5 port map( clk => clk, rst => rst, 
                           req(5) => rq_vc_out(5), req(4) => rq_vc_out(4), 
                           req(3) => rq_vc_out(3), req(2) => rq_vc_out(2), 
                           req(1) => rq_vc_out(1), req(0) => rq_vc_out(0), ack 
                           => vc_available, grant(5) => grant_5_port, grant(4) 
                           => grant_4_port, grant(3) => grant_3_port, grant(2) 
                           => grant_2_port, grant(1) => grant_1_port, grant(0) 
                           => grant_0_port);
   vc_sel_enc_int_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n10, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           vc_sel_enc_1_0_port);
   crossbar_sels_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n12, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_5_port);
   crossbar_sels_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n11, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_4_port);
   vc_sel_enc_int_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n9, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           vc_sel_enc_0_0_port);
   crossbar_sels_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n15, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_2_port);
   crossbar_sels_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n14, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_1_port);
   crossbar_sels_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK
                           => clk, RESET => n8, SET => n5, QN => n124);
   crossbar_sels_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n3, CLK
                           => clk, RESET => n8, SET => n5, QN => n125);
   output_vc_in_use_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2
                           , CLK => clk, RESET => n8, SET => n5, QN => 
                           output_vc_in_use_0_port);
   output_vc_in_use_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1
                           , CLK => clk, RESET => n8, SET => n5, QN => 
                           output_vc_in_use_1_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n5);
   U4 : OA21x2_ASAP7_75t_R port map( A1 => n95, A2 => n94, B => n13, Y => n1);
   U5 : AOI21xp5_ASAP7_75t_R port map( A1 => n118, A2 => n117, B => n119, Y => 
                           n2);
   U6 : AOI22xp5_ASAP7_75t_R port map( A1 => n17, A2 => n119, B1 => n16, B2 => 
                           crossbar_ctrl_vec_0_port, Y => n3);
   U7 : AOI22xp5_ASAP7_75t_R port map( A1 => n17, A2 => n122, B1 => n13, B2 => 
                           crossbar_ctrl_vec_3_port, Y => n4);
   U8 : NOR4xp25_ASAP7_75t_R port map( A => n17, B => grant_0_port, C => 
                           grant_2_port, D => grant_4_port, Y => n103);
   U9 : NOR3xp33_ASAP7_75t_R port map( A => grant_3_port, B => grant_5_port, C 
                           => grant_1_port, Y => n99);
   U10 : NOR2xp33_ASAP7_75t_R port map( A => grant_5_port, B => grant_4_port, Y
                           => n121);
   U11 : NOR2xp33_ASAP7_75t_R port map( A => grant_3_port, B => grant_2_port, Y
                           => n123);
   U12 : INVx1_ASAP7_75t_R port map( A => rst, Y => n8);
   U13 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n21
                           , Y => n91);
   U14 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n20
                           , Y => n82);
   U15 : NOR3xp33_ASAP7_75t_R port map( A => n113, B => 
                           crossbar_ctrl_vec_2_port, C => 
                           crossbar_ctrl_vec_1_port, Y => n114);
   U16 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_0_port, B => n31
                           , Y => n112);
   U17 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n22
                           , Y => n39);
   U18 : HB1xp67_ASAP7_75t_R port map( A => n124, Y => crossbar_ctrl_vec_3_port
                           );
   U19 : HB1xp67_ASAP7_75t_R port map( A => n125, Y => crossbar_ctrl_vec_0_port
                           );
   U20 : NOR2xp33_ASAP7_75t_R port map( A => n103, B => output_vc_in_use_0_port
                           , Y => n119);
   U21 : NOR3xp33_ASAP7_75t_R port map( A => n103, B => output_vc_in_use_1_port
                           , C => n26, Y => n122);
   U22 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n32
                           , Y => n90);
   U29 : INVx1_ASAP7_75t_R port map( A => n33, Y => n9);
   U32 : INVx1_ASAP7_75t_R port map( A => n36, Y => n10);
   U43 : INVx1_ASAP7_75t_R port map( A => n38, Y => n11);
   U44 : INVx1_ASAP7_75t_R port map( A => n37, Y => n12);
   U45 : INVx1_ASAP7_75t_R port map( A => n122, Y => n13);
   U46 : INVx1_ASAP7_75t_R port map( A => n35, Y => n14);
   U47 : INVx1_ASAP7_75t_R port map( A => n34, Y => n15);
   U48 : INVx1_ASAP7_75t_R port map( A => n119, Y => n16);
   U49 : INVx1_ASAP7_75t_R port map( A => n99, Y => n17);
   U50 : INVx1_ASAP7_75t_R port map( A => n121, Y => n18);
   U51 : INVx1_ASAP7_75t_R port map( A => n123, Y => n19);
   U56 : INVx1_ASAP7_75t_R port map( A => packet_end(4), Y => n20);
   U57 : INVx1_ASAP7_75t_R port map( A => packet_end(5), Y => n21);
   U59 : INVx1_ASAP7_75t_R port map( A => packet_end(8), Y => n22);
   U60 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_1_port, Y => n23);
   U61 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_2_port, Y => n24);
   U62 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_0_0_port, Y => n25);
   U63 : INVx1_ASAP7_75t_R port map( A => output_vc_in_use_0_port, Y => n26);
   U64 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_4_port, Y => n27);
   U65 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_5_port, Y => n28);
   U66 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_1_0_port, Y => n29);
   U67 : INVx1_ASAP7_75t_R port map( A => packet_end(0), Y => n30);
   U68 : INVx1_ASAP7_75t_R port map( A => packet_end(1), Y => n31);
   U69 : INVx1_ASAP7_75t_R port map( A => packet_end(9), Y => n32);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity vc_output_allocator_port_num7_vc_num_out2_4 is

   port( clk, rst : in std_logic;  rq_vc_out : in std_logic_vector (5 downto 0)
         ;  granted_vc, packet_end : in std_logic_vector (11 downto 0);  
         crossbar_ctrl_vec : out std_logic_vector (5 downto 0);  vc_sel_enc, 
         output_vc_in_use : out std_logic_vector (1 downto 0);  ack_rq_vc_out :
         out std_logic_vector (5 downto 0));

end vc_output_allocator_port_num7_vc_num_out2_4;

architecture SYN_rtl of vc_output_allocator_port_num7_vc_num_out2_4 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component rr_arbiter_no_delay_CNT6_4
      port( clk, rst : in std_logic;  req : in std_logic_vector (5 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (5 downto 0));
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI211xp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OA211x2_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1O1Ixp25_ASAP7_75t_R
      port( A1, A2, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal crossbar_ctrl_vec_5_port, crossbar_ctrl_vec_4_port, n124, 
      crossbar_ctrl_vec_2_port, crossbar_ctrl_vec_1_port, n125, 
      vc_sel_enc_1_0_port, vc_sel_enc_0_0_port, output_vc_in_use_1_port, 
      output_vc_in_use_0_port, vc_available, grant_5_port, grant_4_port, 
      grant_3_port, grant_2_port, grant_1_port, grant_0_port, n1, n2, n3, n4, 
      n5, crossbar_ctrl_vec_3_port, crossbar_ctrl_vec_0_port, n8, n9, n10, n11,
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123 : std_logic;

begin
   crossbar_ctrl_vec <= ( crossbar_ctrl_vec_5_port, crossbar_ctrl_vec_4_port, 
      crossbar_ctrl_vec_3_port, crossbar_ctrl_vec_2_port, 
      crossbar_ctrl_vec_1_port, crossbar_ctrl_vec_0_port );
   vc_sel_enc <= ( vc_sel_enc_1_0_port, vc_sel_enc_0_0_port );
   output_vc_in_use <= ( output_vc_in_use_1_port, output_vc_in_use_0_port );
   
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => n123, A2 => n13, B1 => n122, B2 
                           => n28, Y => n38);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => n121, A2 => n13, B1 => n122, B2 
                           => n29, Y => n37);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => n120, A2 => n13, B1 => n122, B2 
                           => n30, Y => n36);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => n123, A2 => n16, B1 => n119, B2 
                           => n24, Y => n35);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => n121, A2 => n16, B1 => n119, B2 
                           => n25, Y => n34);
   U28 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n116, A2 => n115, B => n26, C 
                           => n114, Y => n117);
   U30 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n23, B => n110, C => vc_sel_enc_0_0_port, Y => n111)
                           ;
   U31 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(2), B => 
                           crossbar_ctrl_vec_0_port, Y => n110);
   U33 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n21, B => n109, C => n25, Y => n115);
   U34 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(10), B => 
                           crossbar_ctrl_vec_0_port, Y => n109);
   U35 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n31, B => n108, C => n24, Y => n116);
   U36 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(6), B => 
                           crossbar_ctrl_vec_0_port, Y => n108);
   U37 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n107, A2 => n106, B => 
                           vc_sel_enc_0_0_port, C => n27, Y => n118);
   U38 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n20, B => n105, C => n25, Y => n106);
   U39 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(11), B => 
                           crossbar_ctrl_vec_0_port, Y => n105);
   U40 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n32, B => n104, C => n24, Y => n107);
   U41 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(7), B => 
                           crossbar_ctrl_vec_0_port, Y => n104);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => n120, A2 => n16, B1 => n119, B2 
                           => n26, Y => n33);
   U52 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_3_port, A2 =>
                           n22, B => n84, C => n30, Y => n85);
   U53 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(3), B => 
                           crossbar_ctrl_vec_3_port, Y => n84);
   U54 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_3_port, A2 =>
                           n23, B => n83, C => vc_sel_enc_1_0_port, Y => n86);
   U55 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(2), B => 
                           crossbar_ctrl_vec_3_port, Y => n83);
   U58 : NAND2xp5_ASAP7_75t_R port map( A => output_vc_in_use_1_port, B => 
                           output_vc_in_use_0_port, Y => vc_available);
   U81 : A2O1A1O1Ixp25_ASAP7_75t_R port map( A1 => packet_end(3), A2 => 
                           crossbar_ctrl_vec_0_port, B => n112, C => 
                           vc_sel_enc_0_0_port, D => n111, Y => n113);
   U82 : OA211x2_ASAP7_75t_R port map( A1 => n19, A2 => n102, B => n101, C => 
                           n100, Y => n120);
   U83 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(9), A2 => n99, B =>
                           n98, C => n18, Y => n100);
   U84 : AND2x2_ASAP7_75t_R port map( A => granted_vc(11), B => n17, Y => n98);
   U85 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(5), A2 => n99, B =>
                           n97, C => n19, Y => n101);
   U86 : AND2x2_ASAP7_75t_R port map( A => granted_vc(7), B => n17, Y => n97);
   U87 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(1), A2 => n99, B =>
                           n96, C => n121, Y => n102);
   U88 : AND2x2_ASAP7_75t_R port map( A => granted_vc(3), B => n17, Y => n96);
   U89 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n93, A2 => n92, B => n30, C =>
                           output_vc_in_use_1_port, Y => n94);
   U90 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(7), A2 => 
                           crossbar_ctrl_vec_3_port, B => n91, C => 
                           crossbar_ctrl_vec_4_port, Y => n92);
   U91 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(11), A2 => 
                           crossbar_ctrl_vec_3_port, B => n90, C => 
                           crossbar_ctrl_vec_5_port, Y => n93);
   U92 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n89, A2 => n88, B => 
                           vc_sel_enc_1_0_port, C => n87, Y => n95);
   U93 : OAI211xp5_ASAP7_75t_R port map( A1 => n86, A2 => n85, B => n28, C => 
                           n29, Y => n87);
   U94 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(6), A2 => 
                           crossbar_ctrl_vec_3_port, B => n82, C => 
                           crossbar_ctrl_vec_4_port, Y => n88);
   U95 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(10), A2 => 
                           crossbar_ctrl_vec_3_port, B => n39, C => 
                           crossbar_ctrl_vec_5_port, Y => n89);
   U96 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_5_port, Y 
                           => ack_rq_vc_out(5));
   U97 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_4_port, Y 
                           => ack_rq_vc_out(4));
   U98 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_3_port, Y 
                           => ack_rq_vc_out(3));
   U99 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_2_port, Y 
                           => ack_rq_vc_out(2));
   U100 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_1_port, Y 
                           => ack_rq_vc_out(1));
   U101 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_0_port, Y 
                           => ack_rq_vc_out(0));
   rr_arbiter : rr_arbiter_no_delay_CNT6_4 port map( clk => clk, rst => rst, 
                           req(5) => rq_vc_out(5), req(4) => rq_vc_out(4), 
                           req(3) => rq_vc_out(3), req(2) => rq_vc_out(2), 
                           req(1) => rq_vc_out(1), req(0) => rq_vc_out(0), ack 
                           => vc_available, grant(5) => grant_5_port, grant(4) 
                           => grant_4_port, grant(3) => grant_3_port, grant(2) 
                           => grant_2_port, grant(1) => grant_1_port, grant(0) 
                           => grant_0_port);
   vc_sel_enc_int_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n10, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           vc_sel_enc_1_0_port);
   crossbar_sels_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n11, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_4_port);
   crossbar_sels_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n12, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_5_port);
   crossbar_sels_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK
                           => clk, RESET => n8, SET => n5, QN => n124);
   vc_sel_enc_int_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n9, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           vc_sel_enc_0_0_port);
   crossbar_sels_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n15, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_2_port);
   crossbar_sels_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n14, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_1_port);
   crossbar_sels_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n3, CLK
                           => clk, RESET => n8, SET => n5, QN => n125);
   output_vc_in_use_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2
                           , CLK => clk, RESET => n8, SET => n5, QN => 
                           output_vc_in_use_1_port);
   output_vc_in_use_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1
                           , CLK => clk, RESET => n8, SET => n5, QN => 
                           output_vc_in_use_0_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n5);
   U4 : AOI21xp5_ASAP7_75t_R port map( A1 => n118, A2 => n117, B => n119, Y => 
                           n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => n95, A2 => n94, B => n13, Y => n2);
   U6 : AOI22xp5_ASAP7_75t_R port map( A1 => n17, A2 => n119, B1 => n16, B2 => 
                           crossbar_ctrl_vec_0_port, Y => n3);
   U7 : AOI22xp5_ASAP7_75t_R port map( A1 => n17, A2 => n122, B1 => n13, B2 => 
                           crossbar_ctrl_vec_3_port, Y => n4);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => grant_3_port, B => grant_5_port, C 
                           => grant_1_port, Y => n99);
   U9 : NOR2xp33_ASAP7_75t_R port map( A => grant_5_port, B => grant_4_port, Y 
                           => n121);
   U10 : NOR4xp25_ASAP7_75t_R port map( A => n17, B => grant_0_port, C => 
                           grant_2_port, D => grant_4_port, Y => n103);
   U11 : NOR2xp33_ASAP7_75t_R port map( A => grant_3_port, B => grant_2_port, Y
                           => n123);
   U12 : INVx1_ASAP7_75t_R port map( A => rst, Y => n8);
   U13 : NOR3xp33_ASAP7_75t_R port map( A => n113, B => 
                           crossbar_ctrl_vec_2_port, C => 
                           crossbar_ctrl_vec_1_port, Y => n114);
   U14 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_0_port, B => n22
                           , Y => n112);
   U15 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n21
                           , Y => n39);
   U16 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n20
                           , Y => n90);
   U17 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n31
                           , Y => n82);
   U18 : HB1xp67_ASAP7_75t_R port map( A => n124, Y => crossbar_ctrl_vec_3_port
                           );
   U19 : HB1xp67_ASAP7_75t_R port map( A => n125, Y => crossbar_ctrl_vec_0_port
                           );
   U20 : NOR2xp33_ASAP7_75t_R port map( A => n103, B => output_vc_in_use_0_port
                           , Y => n119);
   U21 : NOR3xp33_ASAP7_75t_R port map( A => n103, B => output_vc_in_use_1_port
                           , C => n27, Y => n122);
   U22 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n32
                           , Y => n91);
   U29 : INVx1_ASAP7_75t_R port map( A => n33, Y => n9);
   U32 : INVx1_ASAP7_75t_R port map( A => n36, Y => n10);
   U43 : INVx1_ASAP7_75t_R port map( A => n38, Y => n11);
   U44 : INVx1_ASAP7_75t_R port map( A => n37, Y => n12);
   U45 : INVx1_ASAP7_75t_R port map( A => n122, Y => n13);
   U46 : INVx1_ASAP7_75t_R port map( A => n35, Y => n14);
   U47 : INVx1_ASAP7_75t_R port map( A => n34, Y => n15);
   U48 : INVx1_ASAP7_75t_R port map( A => n119, Y => n16);
   U49 : INVx1_ASAP7_75t_R port map( A => n99, Y => n17);
   U50 : INVx1_ASAP7_75t_R port map( A => n121, Y => n18);
   U51 : INVx1_ASAP7_75t_R port map( A => n123, Y => n19);
   U56 : INVx1_ASAP7_75t_R port map( A => packet_end(9), Y => n20);
   U57 : INVx1_ASAP7_75t_R port map( A => packet_end(8), Y => n21);
   U59 : INVx1_ASAP7_75t_R port map( A => packet_end(1), Y => n22);
   U60 : INVx1_ASAP7_75t_R port map( A => packet_end(0), Y => n23);
   U61 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_1_port, Y => n24);
   U62 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_2_port, Y => n25);
   U63 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_0_0_port, Y => n26);
   U64 : INVx1_ASAP7_75t_R port map( A => output_vc_in_use_0_port, Y => n27);
   U65 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_4_port, Y => n28);
   U66 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_5_port, Y => n29);
   U67 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_1_0_port, Y => n30);
   U68 : INVx1_ASAP7_75t_R port map( A => packet_end(4), Y => n31);
   U69 : INVx1_ASAP7_75t_R port map( A => packet_end(5), Y => n32);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity vc_output_allocator_port_num7_vc_num_out2_3 is

   port( clk, rst : in std_logic;  rq_vc_out : in std_logic_vector (5 downto 0)
         ;  granted_vc, packet_end : in std_logic_vector (11 downto 0);  
         crossbar_ctrl_vec : out std_logic_vector (5 downto 0);  vc_sel_enc, 
         output_vc_in_use : out std_logic_vector (1 downto 0);  ack_rq_vc_out :
         out std_logic_vector (5 downto 0));

end vc_output_allocator_port_num7_vc_num_out2_3;

architecture SYN_rtl of vc_output_allocator_port_num7_vc_num_out2_3 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component rr_arbiter_no_delay_CNT6_3
      port( clk, rst : in std_logic;  req : in std_logic_vector (5 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (5 downto 0));
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI211xp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OA211x2_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1O1Ixp25_ASAP7_75t_R
      port( A1, A2, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal crossbar_ctrl_vec_5_port, crossbar_ctrl_vec_4_port, n124, 
      crossbar_ctrl_vec_2_port, crossbar_ctrl_vec_1_port, n125, 
      vc_sel_enc_1_0_port, vc_sel_enc_0_0_port, output_vc_in_use_1_port, 
      output_vc_in_use_0_port, vc_available, grant_5_port, grant_4_port, 
      grant_3_port, grant_2_port, grant_1_port, grant_0_port, n1, n2, n3, n4, 
      n5, crossbar_ctrl_vec_3_port, crossbar_ctrl_vec_0_port, n8, n9, n10, n11,
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123 : std_logic;

begin
   crossbar_ctrl_vec <= ( crossbar_ctrl_vec_5_port, crossbar_ctrl_vec_4_port, 
      crossbar_ctrl_vec_3_port, crossbar_ctrl_vec_2_port, 
      crossbar_ctrl_vec_1_port, crossbar_ctrl_vec_0_port );
   vc_sel_enc <= ( vc_sel_enc_1_0_port, vc_sel_enc_0_0_port );
   output_vc_in_use <= ( output_vc_in_use_1_port, output_vc_in_use_0_port );
   
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => n123, A2 => n13, B1 => n122, B2 
                           => n29, Y => n38);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => n121, A2 => n13, B1 => n122, B2 
                           => n30, Y => n37);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => n120, A2 => n13, B1 => n122, B2 
                           => n31, Y => n36);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => n123, A2 => n16, B1 => n119, B2 
                           => n25, Y => n35);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => n121, A2 => n16, B1 => n119, B2 
                           => n26, Y => n34);
   U28 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n116, A2 => n115, B => n27, C 
                           => n114, Y => n117);
   U30 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n20, B => n110, C => vc_sel_enc_0_0_port, Y => n111)
                           ;
   U31 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(2), B => 
                           crossbar_ctrl_vec_0_port, Y => n110);
   U33 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n24, B => n109, C => n26, Y => n115);
   U34 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(10), B => 
                           crossbar_ctrl_vec_0_port, Y => n109);
   U35 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n22, B => n108, C => n25, Y => n116);
   U36 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(6), B => 
                           crossbar_ctrl_vec_0_port, Y => n108);
   U37 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n107, A2 => n106, B => 
                           vc_sel_enc_0_0_port, C => n28, Y => n118);
   U38 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n23, B => n105, C => n26, Y => n106);
   U39 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(11), B => 
                           crossbar_ctrl_vec_0_port, Y => n105);
   U40 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n32, B => n104, C => n25, Y => n107);
   U41 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(7), B => 
                           crossbar_ctrl_vec_0_port, Y => n104);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => n120, A2 => n16, B1 => n119, B2 
                           => n27, Y => n33);
   U52 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_3_port, A2 =>
                           n21, B => n84, C => n31, Y => n85);
   U53 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(3), B => 
                           crossbar_ctrl_vec_3_port, Y => n84);
   U54 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_3_port, A2 =>
                           n20, B => n83, C => vc_sel_enc_1_0_port, Y => n86);
   U55 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(2), B => 
                           crossbar_ctrl_vec_3_port, Y => n83);
   U58 : NAND2xp5_ASAP7_75t_R port map( A => output_vc_in_use_1_port, B => 
                           output_vc_in_use_0_port, Y => vc_available);
   U81 : A2O1A1O1Ixp25_ASAP7_75t_R port map( A1 => packet_end(3), A2 => 
                           crossbar_ctrl_vec_0_port, B => n112, C => 
                           vc_sel_enc_0_0_port, D => n111, Y => n113);
   U82 : OA211x2_ASAP7_75t_R port map( A1 => n19, A2 => n102, B => n101, C => 
                           n100, Y => n120);
   U83 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(9), A2 => n99, B =>
                           n98, C => n18, Y => n100);
   U84 : AND2x2_ASAP7_75t_R port map( A => granted_vc(11), B => n17, Y => n98);
   U85 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(5), A2 => n99, B =>
                           n97, C => n19, Y => n101);
   U86 : AND2x2_ASAP7_75t_R port map( A => granted_vc(7), B => n17, Y => n97);
   U87 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(1), A2 => n99, B =>
                           n96, C => n121, Y => n102);
   U88 : AND2x2_ASAP7_75t_R port map( A => granted_vc(3), B => n17, Y => n96);
   U89 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n93, A2 => n92, B => n31, C =>
                           output_vc_in_use_1_port, Y => n94);
   U90 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(7), A2 => 
                           crossbar_ctrl_vec_3_port, B => n91, C => 
                           crossbar_ctrl_vec_4_port, Y => n92);
   U91 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(11), A2 => 
                           crossbar_ctrl_vec_3_port, B => n90, C => 
                           crossbar_ctrl_vec_5_port, Y => n93);
   U92 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n89, A2 => n88, B => 
                           vc_sel_enc_1_0_port, C => n87, Y => n95);
   U93 : OAI211xp5_ASAP7_75t_R port map( A1 => n86, A2 => n85, B => n29, C => 
                           n30, Y => n87);
   U94 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(6), A2 => 
                           crossbar_ctrl_vec_3_port, B => n82, C => 
                           crossbar_ctrl_vec_4_port, Y => n88);
   U95 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(10), A2 => 
                           crossbar_ctrl_vec_3_port, B => n39, C => 
                           crossbar_ctrl_vec_5_port, Y => n89);
   U96 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_5_port, Y 
                           => ack_rq_vc_out(5));
   U97 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_4_port, Y 
                           => ack_rq_vc_out(4));
   U98 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_3_port, Y 
                           => ack_rq_vc_out(3));
   U99 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_2_port, Y 
                           => ack_rq_vc_out(2));
   U100 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_1_port, Y 
                           => ack_rq_vc_out(1));
   U101 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_0_port, Y 
                           => ack_rq_vc_out(0));
   rr_arbiter : rr_arbiter_no_delay_CNT6_3 port map( clk => clk, rst => rst, 
                           req(5) => rq_vc_out(5), req(4) => rq_vc_out(4), 
                           req(3) => rq_vc_out(3), req(2) => rq_vc_out(2), 
                           req(1) => rq_vc_out(1), req(0) => rq_vc_out(0), ack 
                           => vc_available, grant(5) => grant_5_port, grant(4) 
                           => grant_4_port, grant(3) => grant_3_port, grant(2) 
                           => grant_2_port, grant(1) => grant_1_port, grant(0) 
                           => grant_0_port);
   crossbar_sels_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n11, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_4_port);
   crossbar_sels_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n12, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_5_port);
   vc_sel_enc_int_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n10, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           vc_sel_enc_1_0_port);
   crossbar_sels_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK
                           => clk, RESET => n8, SET => n5, QN => n124);
   vc_sel_enc_int_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n9, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           vc_sel_enc_0_0_port);
   crossbar_sels_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n15, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_2_port);
   crossbar_sels_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n14, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_1_port);
   crossbar_sels_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n3, CLK
                           => clk, RESET => n8, SET => n5, QN => n125);
   output_vc_in_use_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2
                           , CLK => clk, RESET => n8, SET => n5, QN => 
                           output_vc_in_use_1_port);
   output_vc_in_use_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1
                           , CLK => clk, RESET => n8, SET => n5, QN => 
                           output_vc_in_use_0_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n5);
   U4 : AOI21xp5_ASAP7_75t_R port map( A1 => n118, A2 => n117, B => n119, Y => 
                           n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => n95, A2 => n94, B => n13, Y => n2);
   U6 : AOI22xp5_ASAP7_75t_R port map( A1 => n17, A2 => n119, B1 => n16, B2 => 
                           crossbar_ctrl_vec_0_port, Y => n3);
   U7 : AOI22xp5_ASAP7_75t_R port map( A1 => n17, A2 => n122, B1 => n13, B2 => 
                           crossbar_ctrl_vec_3_port, Y => n4);
   U8 : NOR4xp25_ASAP7_75t_R port map( A => n17, B => grant_0_port, C => 
                           grant_2_port, D => grant_4_port, Y => n103);
   U9 : NOR2xp33_ASAP7_75t_R port map( A => grant_5_port, B => grant_4_port, Y 
                           => n121);
   U10 : NOR2xp33_ASAP7_75t_R port map( A => grant_3_port, B => grant_2_port, Y
                           => n123);
   U11 : NOR3xp33_ASAP7_75t_R port map( A => grant_3_port, B => grant_5_port, C
                           => grant_1_port, Y => n99);
   U12 : INVx1_ASAP7_75t_R port map( A => rst, Y => n8);
   U13 : NOR3xp33_ASAP7_75t_R port map( A => n113, B => 
                           crossbar_ctrl_vec_2_port, C => 
                           crossbar_ctrl_vec_1_port, Y => n114);
   U14 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_0_port, B => n21
                           , Y => n112);
   U15 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n24
                           , Y => n39);
   U16 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n23
                           , Y => n90);
   U17 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n22
                           , Y => n82);
   U18 : HB1xp67_ASAP7_75t_R port map( A => n124, Y => crossbar_ctrl_vec_3_port
                           );
   U19 : HB1xp67_ASAP7_75t_R port map( A => n125, Y => crossbar_ctrl_vec_0_port
                           );
   U20 : NOR2xp33_ASAP7_75t_R port map( A => n103, B => output_vc_in_use_0_port
                           , Y => n119);
   U21 : NOR3xp33_ASAP7_75t_R port map( A => n103, B => output_vc_in_use_1_port
                           , C => n28, Y => n122);
   U22 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n32
                           , Y => n91);
   U29 : INVx1_ASAP7_75t_R port map( A => n33, Y => n9);
   U32 : INVx1_ASAP7_75t_R port map( A => n36, Y => n10);
   U43 : INVx1_ASAP7_75t_R port map( A => n38, Y => n11);
   U44 : INVx1_ASAP7_75t_R port map( A => n37, Y => n12);
   U45 : INVx1_ASAP7_75t_R port map( A => n122, Y => n13);
   U46 : INVx1_ASAP7_75t_R port map( A => n35, Y => n14);
   U47 : INVx1_ASAP7_75t_R port map( A => n34, Y => n15);
   U48 : INVx1_ASAP7_75t_R port map( A => n119, Y => n16);
   U49 : INVx1_ASAP7_75t_R port map( A => n99, Y => n17);
   U50 : INVx1_ASAP7_75t_R port map( A => n121, Y => n18);
   U51 : INVx1_ASAP7_75t_R port map( A => n123, Y => n19);
   U56 : INVx1_ASAP7_75t_R port map( A => packet_end(0), Y => n20);
   U57 : INVx1_ASAP7_75t_R port map( A => packet_end(1), Y => n21);
   U59 : INVx1_ASAP7_75t_R port map( A => packet_end(4), Y => n22);
   U60 : INVx1_ASAP7_75t_R port map( A => packet_end(9), Y => n23);
   U61 : INVx1_ASAP7_75t_R port map( A => packet_end(8), Y => n24);
   U62 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_1_port, Y => n25);
   U63 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_2_port, Y => n26);
   U64 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_0_0_port, Y => n27);
   U65 : INVx1_ASAP7_75t_R port map( A => output_vc_in_use_0_port, Y => n28);
   U66 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_4_port, Y => n29);
   U67 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_5_port, Y => n30);
   U68 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_1_0_port, Y => n31);
   U69 : INVx1_ASAP7_75t_R port map( A => packet_end(5), Y => n32);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity vc_output_allocator_port_num7_vc_num_out2_2 is

   port( clk, rst : in std_logic;  rq_vc_out : in std_logic_vector (5 downto 0)
         ;  granted_vc, packet_end : in std_logic_vector (11 downto 0);  
         crossbar_ctrl_vec : out std_logic_vector (5 downto 0);  vc_sel_enc, 
         output_vc_in_use : out std_logic_vector (1 downto 0);  ack_rq_vc_out :
         out std_logic_vector (5 downto 0));

end vc_output_allocator_port_num7_vc_num_out2_2;

architecture SYN_rtl of vc_output_allocator_port_num7_vc_num_out2_2 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component rr_arbiter_no_delay_CNT6_2
      port( clk, rst : in std_logic;  req : in std_logic_vector (5 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (5 downto 0));
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI211xp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OA211x2_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1O1Ixp25_ASAP7_75t_R
      port( A1, A2, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal crossbar_ctrl_vec_5_port, crossbar_ctrl_vec_4_port, n124, 
      crossbar_ctrl_vec_2_port, crossbar_ctrl_vec_1_port, n125, 
      vc_sel_enc_1_0_port, vc_sel_enc_0_0_port, output_vc_in_use_1_port, 
      output_vc_in_use_0_port, vc_available, grant_5_port, grant_4_port, 
      grant_3_port, grant_2_port, grant_1_port, grant_0_port, n1, n2, n3, n4, 
      n5, crossbar_ctrl_vec_3_port, crossbar_ctrl_vec_0_port, n8, n9, n10, n11,
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123 : std_logic;

begin
   crossbar_ctrl_vec <= ( crossbar_ctrl_vec_5_port, crossbar_ctrl_vec_4_port, 
      crossbar_ctrl_vec_3_port, crossbar_ctrl_vec_2_port, 
      crossbar_ctrl_vec_1_port, crossbar_ctrl_vec_0_port );
   vc_sel_enc <= ( vc_sel_enc_1_0_port, vc_sel_enc_0_0_port );
   output_vc_in_use <= ( output_vc_in_use_1_port, output_vc_in_use_0_port );
   
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => n123, A2 => n13, B1 => n122, B2 
                           => n30, Y => n38);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => n121, A2 => n13, B1 => n122, B2 
                           => n31, Y => n37);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => n120, A2 => n13, B1 => n122, B2 
                           => n32, Y => n36);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => n123, A2 => n16, B1 => n119, B2 
                           => n26, Y => n35);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => n121, A2 => n16, B1 => n119, B2 
                           => n27, Y => n34);
   U28 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n116, A2 => n115, B => n28, C 
                           => n114, Y => n117);
   U30 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n23, B => n110, C => vc_sel_enc_0_0_port, Y => n111)
                           ;
   U31 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(2), B => 
                           crossbar_ctrl_vec_0_port, Y => n110);
   U33 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n25, B => n109, C => n27, Y => n115);
   U34 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(10), B => 
                           crossbar_ctrl_vec_0_port, Y => n109);
   U35 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n21, B => n108, C => n26, Y => n116);
   U36 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(6), B => 
                           crossbar_ctrl_vec_0_port, Y => n108);
   U37 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n107, A2 => n106, B => 
                           vc_sel_enc_0_0_port, C => n29, Y => n118);
   U38 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n24, B => n105, C => n27, Y => n106);
   U39 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(11), B => 
                           crossbar_ctrl_vec_0_port, Y => n105);
   U40 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n20, B => n104, C => n26, Y => n107);
   U41 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(7), B => 
                           crossbar_ctrl_vec_0_port, Y => n104);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => n120, A2 => n16, B1 => n119, B2 
                           => n28, Y => n33);
   U52 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_3_port, A2 =>
                           n22, B => n84, C => n32, Y => n85);
   U53 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(3), B => 
                           crossbar_ctrl_vec_3_port, Y => n84);
   U54 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_3_port, A2 =>
                           n23, B => n83, C => vc_sel_enc_1_0_port, Y => n86);
   U55 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(2), B => 
                           crossbar_ctrl_vec_3_port, Y => n83);
   U58 : NAND2xp5_ASAP7_75t_R port map( A => output_vc_in_use_1_port, B => 
                           output_vc_in_use_0_port, Y => vc_available);
   U81 : A2O1A1O1Ixp25_ASAP7_75t_R port map( A1 => packet_end(3), A2 => 
                           crossbar_ctrl_vec_0_port, B => n112, C => 
                           vc_sel_enc_0_0_port, D => n111, Y => n113);
   U82 : OA211x2_ASAP7_75t_R port map( A1 => n19, A2 => n102, B => n101, C => 
                           n100, Y => n120);
   U83 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(9), A2 => n99, B =>
                           n98, C => n18, Y => n100);
   U84 : AND2x2_ASAP7_75t_R port map( A => granted_vc(11), B => n17, Y => n98);
   U85 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(5), A2 => n99, B =>
                           n97, C => n19, Y => n101);
   U86 : AND2x2_ASAP7_75t_R port map( A => granted_vc(7), B => n17, Y => n97);
   U87 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(1), A2 => n99, B =>
                           n96, C => n121, Y => n102);
   U88 : AND2x2_ASAP7_75t_R port map( A => granted_vc(3), B => n17, Y => n96);
   U89 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n93, A2 => n92, B => n32, C =>
                           output_vc_in_use_1_port, Y => n94);
   U90 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(7), A2 => 
                           crossbar_ctrl_vec_3_port, B => n91, C => 
                           crossbar_ctrl_vec_4_port, Y => n92);
   U91 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(11), A2 => 
                           crossbar_ctrl_vec_3_port, B => n90, C => 
                           crossbar_ctrl_vec_5_port, Y => n93);
   U92 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n89, A2 => n88, B => 
                           vc_sel_enc_1_0_port, C => n87, Y => n95);
   U93 : OAI211xp5_ASAP7_75t_R port map( A1 => n86, A2 => n85, B => n30, C => 
                           n31, Y => n87);
   U94 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(6), A2 => 
                           crossbar_ctrl_vec_3_port, B => n82, C => 
                           crossbar_ctrl_vec_4_port, Y => n88);
   U95 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(10), A2 => 
                           crossbar_ctrl_vec_3_port, B => n39, C => 
                           crossbar_ctrl_vec_5_port, Y => n89);
   U96 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_5_port, Y 
                           => ack_rq_vc_out(5));
   U97 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_4_port, Y 
                           => ack_rq_vc_out(4));
   U98 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_3_port, Y 
                           => ack_rq_vc_out(3));
   U99 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_2_port, Y 
                           => ack_rq_vc_out(2));
   U100 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_1_port, Y 
                           => ack_rq_vc_out(1));
   U101 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_0_port, Y 
                           => ack_rq_vc_out(0));
   rr_arbiter : rr_arbiter_no_delay_CNT6_2 port map( clk => clk, rst => rst, 
                           req(5) => rq_vc_out(5), req(4) => rq_vc_out(4), 
                           req(3) => rq_vc_out(3), req(2) => rq_vc_out(2), 
                           req(1) => rq_vc_out(1), req(0) => rq_vc_out(0), ack 
                           => vc_available, grant(5) => grant_5_port, grant(4) 
                           => grant_4_port, grant(3) => grant_3_port, grant(2) 
                           => grant_2_port, grant(1) => grant_1_port, grant(0) 
                           => grant_0_port);
   vc_sel_enc_int_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n10, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           vc_sel_enc_1_0_port);
   crossbar_sels_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n11, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_4_port);
   crossbar_sels_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n12, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_5_port);
   crossbar_sels_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK
                           => clk, RESET => n8, SET => n5, QN => n124);
   vc_sel_enc_int_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n9, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           vc_sel_enc_0_0_port);
   crossbar_sels_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n15, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_2_port);
   crossbar_sels_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n14, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_1_port);
   crossbar_sels_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n3, CLK
                           => clk, RESET => n8, SET => n5, QN => n125);
   output_vc_in_use_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2
                           , CLK => clk, RESET => n8, SET => n5, QN => 
                           output_vc_in_use_1_port);
   output_vc_in_use_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1
                           , CLK => clk, RESET => n8, SET => n5, QN => 
                           output_vc_in_use_0_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n5);
   U4 : AOI21xp5_ASAP7_75t_R port map( A1 => n118, A2 => n117, B => n119, Y => 
                           n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => n95, A2 => n94, B => n13, Y => n2);
   U6 : AOI22xp5_ASAP7_75t_R port map( A1 => n17, A2 => n119, B1 => n16, B2 => 
                           crossbar_ctrl_vec_0_port, Y => n3);
   U7 : AOI22xp5_ASAP7_75t_R port map( A1 => n17, A2 => n122, B1 => n13, B2 => 
                           crossbar_ctrl_vec_3_port, Y => n4);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => grant_3_port, B => grant_5_port, C 
                           => grant_1_port, Y => n99);
   U9 : NOR4xp25_ASAP7_75t_R port map( A => n17, B => grant_0_port, C => 
                           grant_2_port, D => grant_4_port, Y => n103);
   U10 : NOR2xp33_ASAP7_75t_R port map( A => grant_5_port, B => grant_4_port, Y
                           => n121);
   U11 : NOR2xp33_ASAP7_75t_R port map( A => grant_3_port, B => grant_2_port, Y
                           => n123);
   U12 : INVx1_ASAP7_75t_R port map( A => rst, Y => n8);
   U13 : NOR3xp33_ASAP7_75t_R port map( A => n113, B => 
                           crossbar_ctrl_vec_2_port, C => 
                           crossbar_ctrl_vec_1_port, Y => n114);
   U14 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_0_port, B => n22
                           , Y => n112);
   U15 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n21
                           , Y => n82);
   U16 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n20
                           , Y => n91);
   U17 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n24
                           , Y => n90);
   U18 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n25
                           , Y => n39);
   U19 : HB1xp67_ASAP7_75t_R port map( A => n124, Y => crossbar_ctrl_vec_3_port
                           );
   U20 : HB1xp67_ASAP7_75t_R port map( A => n125, Y => crossbar_ctrl_vec_0_port
                           );
   U21 : NOR2xp33_ASAP7_75t_R port map( A => n103, B => output_vc_in_use_0_port
                           , Y => n119);
   U22 : NOR3xp33_ASAP7_75t_R port map( A => n103, B => output_vc_in_use_1_port
                           , C => n29, Y => n122);
   U29 : INVx1_ASAP7_75t_R port map( A => n33, Y => n9);
   U32 : INVx1_ASAP7_75t_R port map( A => n36, Y => n10);
   U43 : INVx1_ASAP7_75t_R port map( A => n38, Y => n11);
   U44 : INVx1_ASAP7_75t_R port map( A => n37, Y => n12);
   U45 : INVx1_ASAP7_75t_R port map( A => n122, Y => n13);
   U46 : INVx1_ASAP7_75t_R port map( A => n35, Y => n14);
   U47 : INVx1_ASAP7_75t_R port map( A => n34, Y => n15);
   U48 : INVx1_ASAP7_75t_R port map( A => n119, Y => n16);
   U49 : INVx1_ASAP7_75t_R port map( A => n99, Y => n17);
   U50 : INVx1_ASAP7_75t_R port map( A => n121, Y => n18);
   U51 : INVx1_ASAP7_75t_R port map( A => n123, Y => n19);
   U56 : INVx1_ASAP7_75t_R port map( A => packet_end(5), Y => n20);
   U57 : INVx1_ASAP7_75t_R port map( A => packet_end(4), Y => n21);
   U59 : INVx1_ASAP7_75t_R port map( A => packet_end(1), Y => n22);
   U60 : INVx1_ASAP7_75t_R port map( A => packet_end(0), Y => n23);
   U61 : INVx1_ASAP7_75t_R port map( A => packet_end(9), Y => n24);
   U62 : INVx1_ASAP7_75t_R port map( A => packet_end(8), Y => n25);
   U63 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_1_port, Y => n26);
   U64 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_2_port, Y => n27);
   U65 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_0_0_port, Y => n28);
   U66 : INVx1_ASAP7_75t_R port map( A => output_vc_in_use_0_port, Y => n29);
   U67 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_4_port, Y => n30);
   U68 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_5_port, Y => n31);
   U69 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_1_0_port, Y => n32);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity vc_output_allocator_port_num7_vc_num_out2_1 is

   port( clk, rst : in std_logic;  rq_vc_out : in std_logic_vector (5 downto 0)
         ;  granted_vc, packet_end : in std_logic_vector (11 downto 0);  
         crossbar_ctrl_vec : out std_logic_vector (5 downto 0);  vc_sel_enc, 
         output_vc_in_use : out std_logic_vector (1 downto 0);  ack_rq_vc_out :
         out std_logic_vector (5 downto 0));

end vc_output_allocator_port_num7_vc_num_out2_1;

architecture SYN_rtl of vc_output_allocator_port_num7_vc_num_out2_1 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component rr_arbiter_no_delay_CNT6_1
      port( clk, rst : in std_logic;  req : in std_logic_vector (5 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (5 downto 0));
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI211xp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OA211x2_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1O1Ixp25_ASAP7_75t_R
      port( A1, A2, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal crossbar_ctrl_vec_5_port, crossbar_ctrl_vec_4_port, n124, 
      crossbar_ctrl_vec_2_port, crossbar_ctrl_vec_1_port, n125, 
      vc_sel_enc_1_0_port, vc_sel_enc_0_0_port, output_vc_in_use_1_port, 
      output_vc_in_use_0_port, vc_available, grant_5_port, grant_4_port, 
      grant_3_port, grant_2_port, grant_1_port, grant_0_port, n1, n2, n3, n4, 
      n5, crossbar_ctrl_vec_3_port, crossbar_ctrl_vec_0_port, n8, n9, n10, n11,
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123 : std_logic;

begin
   crossbar_ctrl_vec <= ( crossbar_ctrl_vec_5_port, crossbar_ctrl_vec_4_port, 
      crossbar_ctrl_vec_3_port, crossbar_ctrl_vec_2_port, 
      crossbar_ctrl_vec_1_port, crossbar_ctrl_vec_0_port );
   vc_sel_enc <= ( vc_sel_enc_1_0_port, vc_sel_enc_0_0_port );
   output_vc_in_use <= ( output_vc_in_use_1_port, output_vc_in_use_0_port );
   
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => n123, A2 => n13, B1 => n122, B2 
                           => n25, Y => n38);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => n121, A2 => n13, B1 => n122, B2 
                           => n26, Y => n37);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => n120, A2 => n13, B1 => n122, B2 
                           => n27, Y => n36);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => n123, A2 => n16, B1 => n119, B2 
                           => n21, Y => n35);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => n121, A2 => n16, B1 => n119, B2 
                           => n22, Y => n34);
   U28 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n116, A2 => n115, B => n23, C 
                           => n114, Y => n117);
   U30 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n20, B => n110, C => vc_sel_enc_0_0_port, Y => n111)
                           ;
   U31 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(2), B => 
                           crossbar_ctrl_vec_0_port, Y => n110);
   U33 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n31, B => n109, C => n22, Y => n115);
   U34 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(10), B => 
                           crossbar_ctrl_vec_0_port, Y => n109);
   U35 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n29, B => n108, C => n21, Y => n116);
   U36 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(6), B => 
                           crossbar_ctrl_vec_0_port, Y => n108);
   U37 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n107, A2 => n106, B => 
                           vc_sel_enc_0_0_port, C => n24, Y => n118);
   U38 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n32, B => n105, C => n22, Y => n106);
   U39 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(11), B => 
                           crossbar_ctrl_vec_0_port, Y => n105);
   U40 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n30, B => n104, C => n21, Y => n107);
   U41 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(7), B => 
                           crossbar_ctrl_vec_0_port, Y => n104);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => n120, A2 => n16, B1 => n119, B2 
                           => n23, Y => n33);
   U52 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_3_port, A2 =>
                           n28, B => n84, C => n27, Y => n85);
   U53 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(3), B => 
                           crossbar_ctrl_vec_3_port, Y => n84);
   U54 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_3_port, A2 =>
                           n20, B => n83, C => vc_sel_enc_1_0_port, Y => n86);
   U55 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(2), B => 
                           crossbar_ctrl_vec_3_port, Y => n83);
   U58 : NAND2xp5_ASAP7_75t_R port map( A => output_vc_in_use_1_port, B => 
                           output_vc_in_use_0_port, Y => vc_available);
   U81 : A2O1A1O1Ixp25_ASAP7_75t_R port map( A1 => packet_end(3), A2 => 
                           crossbar_ctrl_vec_0_port, B => n112, C => 
                           vc_sel_enc_0_0_port, D => n111, Y => n113);
   U82 : OA211x2_ASAP7_75t_R port map( A1 => n19, A2 => n102, B => n101, C => 
                           n100, Y => n120);
   U83 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(9), A2 => n99, B =>
                           n98, C => n18, Y => n100);
   U84 : AND2x2_ASAP7_75t_R port map( A => granted_vc(11), B => n17, Y => n98);
   U85 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(5), A2 => n99, B =>
                           n97, C => n19, Y => n101);
   U86 : AND2x2_ASAP7_75t_R port map( A => granted_vc(7), B => n17, Y => n97);
   U87 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(1), A2 => n99, B =>
                           n96, C => n121, Y => n102);
   U88 : AND2x2_ASAP7_75t_R port map( A => granted_vc(3), B => n17, Y => n96);
   U89 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n93, A2 => n92, B => n27, C =>
                           output_vc_in_use_1_port, Y => n94);
   U90 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(7), A2 => 
                           crossbar_ctrl_vec_3_port, B => n91, C => 
                           crossbar_ctrl_vec_4_port, Y => n92);
   U91 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(11), A2 => 
                           crossbar_ctrl_vec_3_port, B => n90, C => 
                           crossbar_ctrl_vec_5_port, Y => n93);
   U92 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n89, A2 => n88, B => 
                           vc_sel_enc_1_0_port, C => n87, Y => n95);
   U93 : OAI211xp5_ASAP7_75t_R port map( A1 => n86, A2 => n85, B => n25, C => 
                           n26, Y => n87);
   U94 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(6), A2 => 
                           crossbar_ctrl_vec_3_port, B => n82, C => 
                           crossbar_ctrl_vec_4_port, Y => n88);
   U95 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(10), A2 => 
                           crossbar_ctrl_vec_3_port, B => n39, C => 
                           crossbar_ctrl_vec_5_port, Y => n89);
   U96 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_5_port, Y 
                           => ack_rq_vc_out(5));
   U97 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_4_port, Y 
                           => ack_rq_vc_out(4));
   U98 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_3_port, Y 
                           => ack_rq_vc_out(3));
   U99 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_2_port, Y 
                           => ack_rq_vc_out(2));
   U100 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_1_port, Y 
                           => ack_rq_vc_out(1));
   U101 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_0_port, Y 
                           => ack_rq_vc_out(0));
   rr_arbiter : rr_arbiter_no_delay_CNT6_1 port map( clk => clk, rst => rst, 
                           req(5) => rq_vc_out(5), req(4) => rq_vc_out(4), 
                           req(3) => rq_vc_out(3), req(2) => rq_vc_out(2), 
                           req(1) => rq_vc_out(1), req(0) => rq_vc_out(0), ack 
                           => vc_available, grant(5) => grant_5_port, grant(4) 
                           => grant_4_port, grant(3) => grant_3_port, grant(2) 
                           => grant_2_port, grant(1) => grant_1_port, grant(0) 
                           => grant_0_port);
   crossbar_sels_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n11, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_4_port);
   vc_sel_enc_int_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n10, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           vc_sel_enc_1_0_port);
   crossbar_sels_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n12, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_5_port);
   crossbar_sels_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK
                           => clk, RESET => n8, SET => n5, QN => n124);
   crossbar_sels_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n14, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_1_port);
   vc_sel_enc_int_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n9, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           vc_sel_enc_0_0_port);
   crossbar_sels_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n15, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_2_port);
   crossbar_sels_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n3, CLK
                           => clk, RESET => n8, SET => n5, QN => n125);
   output_vc_in_use_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2
                           , CLK => clk, RESET => n8, SET => n5, QN => 
                           output_vc_in_use_1_port);
   output_vc_in_use_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1
                           , CLK => clk, RESET => n8, SET => n5, QN => 
                           output_vc_in_use_0_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n5);
   U4 : AOI21xp5_ASAP7_75t_R port map( A1 => n118, A2 => n117, B => n119, Y => 
                           n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => n95, A2 => n94, B => n13, Y => n2);
   U6 : AOI22xp5_ASAP7_75t_R port map( A1 => n17, A2 => n119, B1 => n16, B2 => 
                           crossbar_ctrl_vec_0_port, Y => n3);
   U7 : AOI22xp5_ASAP7_75t_R port map( A1 => n17, A2 => n122, B1 => n13, B2 => 
                           crossbar_ctrl_vec_3_port, Y => n4);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => grant_3_port, B => grant_5_port, C 
                           => grant_1_port, Y => n99);
   U9 : NOR4xp25_ASAP7_75t_R port map( A => n17, B => grant_0_port, C => 
                           grant_2_port, D => grant_4_port, Y => n103);
   U10 : NOR2xp33_ASAP7_75t_R port map( A => grant_5_port, B => grant_4_port, Y
                           => n121);
   U11 : INVx1_ASAP7_75t_R port map( A => rst, Y => n8);
   U12 : NOR2xp33_ASAP7_75t_R port map( A => grant_3_port, B => grant_2_port, Y
                           => n123);
   U13 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n32
                           , Y => n90);
   U14 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n31
                           , Y => n39);
   U15 : NOR3xp33_ASAP7_75t_R port map( A => n113, B => 
                           crossbar_ctrl_vec_2_port, C => 
                           crossbar_ctrl_vec_1_port, Y => n114);
   U16 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_0_port, B => n28
                           , Y => n112);
   U17 : HB1xp67_ASAP7_75t_R port map( A => n124, Y => crossbar_ctrl_vec_3_port
                           );
   U18 : HB1xp67_ASAP7_75t_R port map( A => n125, Y => crossbar_ctrl_vec_0_port
                           );
   U19 : NOR2xp33_ASAP7_75t_R port map( A => n103, B => output_vc_in_use_0_port
                           , Y => n119);
   U20 : NOR3xp33_ASAP7_75t_R port map( A => n103, B => output_vc_in_use_1_port
                           , C => n24, Y => n122);
   U21 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n30
                           , Y => n91);
   U22 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n29
                           , Y => n82);
   U29 : INVx1_ASAP7_75t_R port map( A => n33, Y => n9);
   U32 : INVx1_ASAP7_75t_R port map( A => n36, Y => n10);
   U43 : INVx1_ASAP7_75t_R port map( A => n38, Y => n11);
   U44 : INVx1_ASAP7_75t_R port map( A => n37, Y => n12);
   U45 : INVx1_ASAP7_75t_R port map( A => n122, Y => n13);
   U46 : INVx1_ASAP7_75t_R port map( A => n35, Y => n14);
   U47 : INVx1_ASAP7_75t_R port map( A => n34, Y => n15);
   U48 : INVx1_ASAP7_75t_R port map( A => n119, Y => n16);
   U49 : INVx1_ASAP7_75t_R port map( A => n99, Y => n17);
   U50 : INVx1_ASAP7_75t_R port map( A => n121, Y => n18);
   U51 : INVx1_ASAP7_75t_R port map( A => n123, Y => n19);
   U56 : INVx1_ASAP7_75t_R port map( A => packet_end(0), Y => n20);
   U57 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_1_port, Y => n21);
   U59 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_2_port, Y => n22);
   U60 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_0_0_port, Y => n23);
   U61 : INVx1_ASAP7_75t_R port map( A => output_vc_in_use_0_port, Y => n24);
   U62 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_4_port, Y => n25);
   U63 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_5_port, Y => n26);
   U64 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_1_0_port, Y => n27);
   U65 : INVx1_ASAP7_75t_R port map( A => packet_end(1), Y => n28);
   U66 : INVx1_ASAP7_75t_R port map( A => packet_end(4), Y => n29);
   U67 : INVx1_ASAP7_75t_R port map( A => packet_end(5), Y => n30);
   U68 : INVx1_ASAP7_75t_R port map( A => packet_end(8), Y => n31);
   U69 : INVx1_ASAP7_75t_R port map( A => packet_end(9), Y => n32);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity fifo_buff_depth2_12 is

   port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, clk, 
         rst : in std_logic;  data_out : out std_logic_vector (63 downto 0);  
         valid_data : out std_logic);

end fifo_buff_depth2_12;

architecture SYN_rtl of fifo_buff_depth2_12 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx3_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal valid_data_port, read_pointer_0_port, fifo_1_63_port, fifo_1_62_port,
      fifo_1_61_port, fifo_1_60_port, fifo_1_59_port, fifo_1_58_port, 
      fifo_1_57_port, fifo_1_56_port, fifo_1_55_port, fifo_1_54_port, 
      fifo_1_53_port, fifo_1_52_port, fifo_1_51_port, fifo_1_50_port, 
      fifo_1_49_port, fifo_1_48_port, fifo_1_47_port, fifo_1_46_port, 
      fifo_1_45_port, fifo_1_44_port, fifo_1_43_port, fifo_1_42_port, 
      fifo_1_41_port, fifo_1_40_port, fifo_1_39_port, fifo_1_38_port, 
      fifo_1_37_port, fifo_1_36_port, fifo_1_35_port, fifo_1_34_port, 
      fifo_1_33_port, fifo_1_32_port, fifo_1_31_port, fifo_1_30_port, 
      fifo_1_29_port, fifo_1_28_port, fifo_1_27_port, fifo_1_26_port, 
      fifo_1_25_port, fifo_1_24_port, fifo_1_23_port, fifo_1_22_port, 
      fifo_1_21_port, fifo_1_20_port, fifo_1_19_port, fifo_1_18_port, 
      fifo_1_17_port, fifo_1_16_port, fifo_1_15_port, fifo_1_14_port, 
      fifo_1_13_port, fifo_1_12_port, fifo_1_11_port, fifo_1_10_port, 
      fifo_1_9_port, fifo_1_8_port, fifo_1_7_port, fifo_1_6_port, fifo_1_5_port
      , fifo_1_4_port, fifo_1_3_port, fifo_1_2_port, fifo_1_1_port, 
      fifo_1_0_port, fifo_0_63_port, fifo_0_62_port, fifo_0_61_port, 
      fifo_0_60_port, fifo_0_59_port, fifo_0_58_port, fifo_0_57_port, 
      fifo_0_56_port, fifo_0_55_port, fifo_0_54_port, fifo_0_53_port, 
      fifo_0_52_port, fifo_0_51_port, fifo_0_50_port, fifo_0_49_port, 
      fifo_0_48_port, fifo_0_47_port, fifo_0_46_port, fifo_0_45_port, 
      fifo_0_44_port, fifo_0_43_port, fifo_0_42_port, fifo_0_41_port, 
      fifo_0_40_port, fifo_0_39_port, fifo_0_38_port, fifo_0_37_port, 
      fifo_0_36_port, fifo_0_35_port, fifo_0_34_port, fifo_0_33_port, 
      fifo_0_32_port, fifo_0_31_port, fifo_0_30_port, fifo_0_29_port, 
      fifo_0_28_port, fifo_0_27_port, fifo_0_26_port, fifo_0_25_port, 
      fifo_0_24_port, fifo_0_23_port, fifo_0_22_port, fifo_0_21_port, 
      fifo_0_20_port, fifo_0_19_port, fifo_0_18_port, fifo_0_17_port, 
      fifo_0_16_port, fifo_0_15_port, fifo_0_14_port, fifo_0_13_port, 
      fifo_0_12_port, fifo_0_11_port, fifo_0_10_port, fifo_0_9_port, 
      fifo_0_8_port, fifo_0_7_port, fifo_0_6_port, fifo_0_5_port, fifo_0_4_port
      , fifo_0_3_port, fifo_0_2_port, fifo_0_1_port, fifo_0_0_port, N7, N9, n1,
      n3, n5, n7_port, n9_port, n11, n13, n15, n17, n19, n21, n23, n25, n27, 
      n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57
      , n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, 
      n87, n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, n111, 
      n113, n115, n117, n119, n121, n123, n125, n127, n129, n131, n133, n135, 
      n137, n139, n141, n143, n145, n147, n149, n151, n153, n155, n157, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238 : std_logic;

begin
   valid_data <= valid_data_port;
   
   U4 : XOR2xp5_ASAP7_75t_R port map( A => N7, B => n43, Y => n238);
   U143 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_9_port, B1 => 
                           n43, B2 => fifo_0_9_port, Y => data_out(9));
   U144 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_8_port, B1 => 
                           n43, B2 => fifo_0_8_port, Y => data_out(8));
   U145 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_7_port, B1 => 
                           n43, B2 => fifo_0_7_port, Y => data_out(7));
   U146 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_6_port, B1 => 
                           n43, B2 => fifo_0_6_port, Y => data_out(6));
   U147 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_63_port, B1 => 
                           n43, B2 => fifo_0_63_port, Y => data_out(63));
   U148 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_62_port, B1 => 
                           n43, B2 => fifo_0_62_port, Y => data_out(62));
   U149 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_61_port, B1 => 
                           n43, B2 => fifo_0_61_port, Y => data_out(61));
   U150 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_60_port, B1 => 
                           n43, B2 => fifo_0_60_port, Y => data_out(60));
   U151 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_5_port, B1 => 
                           n43, B2 => fifo_0_5_port, Y => data_out(5));
   U152 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_59_port, B1 => 
                           n43, B2 => fifo_0_59_port, Y => data_out(59));
   U153 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_58_port, B1 => 
                           n43, B2 => fifo_0_58_port, Y => data_out(58));
   U154 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_57_port, B1 => 
                           n43, B2 => fifo_0_57_port, Y => data_out(57));
   U155 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_56_port, B1 => 
                           n43, B2 => fifo_0_56_port, Y => data_out(56));
   U156 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_55_port, B1 => 
                           n43, B2 => fifo_0_55_port, Y => data_out(55));
   U157 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_54_port, B1 => 
                           n43, B2 => fifo_0_54_port, Y => data_out(54));
   U158 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_53_port, B1 => 
                           n43, B2 => fifo_0_53_port, Y => data_out(53));
   U159 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_52_port, B1 => 
                           n43, B2 => fifo_0_52_port, Y => data_out(52));
   U160 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_51_port, B1 => 
                           n43, B2 => fifo_0_51_port, Y => data_out(51));
   U161 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_50_port, B1 => 
                           n43, B2 => fifo_0_50_port, Y => data_out(50));
   U162 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_4_port, B1 => 
                           n43, B2 => fifo_0_4_port, Y => data_out(4));
   U163 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_49_port, B1 => 
                           n43, B2 => fifo_0_49_port, Y => data_out(49));
   U164 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_48_port, B1 => 
                           n43, B2 => fifo_0_48_port, Y => data_out(48));
   U165 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_47_port, B1 => 
                           n43, B2 => fifo_0_47_port, Y => data_out(47));
   U166 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_46_port, B1 => 
                           n43, B2 => fifo_0_46_port, Y => data_out(46));
   U167 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_45_port, B1 => 
                           n43, B2 => fifo_0_45_port, Y => data_out(45));
   U168 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_44_port, B1 => 
                           n43, B2 => fifo_0_44_port, Y => data_out(44));
   U169 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_43_port, B1 => 
                           n43, B2 => fifo_0_43_port, Y => data_out(43));
   U170 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_42_port, B1 => 
                           n43, B2 => fifo_0_42_port, Y => data_out(42));
   U171 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_41_port, B1 => 
                           n43, B2 => fifo_0_41_port, Y => data_out(41));
   U172 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_40_port, B1 => 
                           n43, B2 => fifo_0_40_port, Y => data_out(40));
   U173 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_3_port, B1 => 
                           n43, B2 => fifo_0_3_port, Y => data_out(3));
   U174 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_39_port, B1 => 
                           n43, B2 => fifo_0_39_port, Y => data_out(39));
   U175 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_38_port, B1 => 
                           n43, B2 => fifo_0_38_port, Y => data_out(38));
   U176 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_37_port, B1 => 
                           n43, B2 => fifo_0_37_port, Y => data_out(37));
   U177 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_36_port, B1 => 
                           n43, B2 => fifo_0_36_port, Y => data_out(36));
   U178 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_35_port, B1 => 
                           n43, B2 => fifo_0_35_port, Y => data_out(35));
   U179 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_34_port, B1 => 
                           n43, B2 => fifo_0_34_port, Y => data_out(34));
   U180 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_33_port, B1 => 
                           n43, B2 => fifo_0_33_port, Y => data_out(33));
   U181 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_32_port, B1 => 
                           n43, B2 => fifo_0_32_port, Y => data_out(32));
   U182 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_31_port, B1 => 
                           n43, B2 => fifo_0_31_port, Y => data_out(31));
   U183 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_30_port, B1 => 
                           n43, B2 => fifo_0_30_port, Y => data_out(30));
   U184 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_2_port, B1 => 
                           n43, B2 => fifo_0_2_port, Y => data_out(2));
   U185 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_29_port, B1 => 
                           n43, B2 => fifo_0_29_port, Y => data_out(29));
   U186 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_28_port, B1 => 
                           n43, B2 => fifo_0_28_port, Y => data_out(28));
   U187 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_27_port, B1 => 
                           n43, B2 => fifo_0_27_port, Y => data_out(27));
   U188 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_26_port, B1 => 
                           n43, B2 => fifo_0_26_port, Y => data_out(26));
   U189 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_25_port, B1 => 
                           n43, B2 => fifo_0_25_port, Y => data_out(25));
   U190 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_24_port, B1 => 
                           n43, B2 => fifo_0_24_port, Y => data_out(24));
   U191 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_23_port, B1 => 
                           n43, B2 => fifo_0_23_port, Y => data_out(23));
   U192 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_22_port, B1 => 
                           n43, B2 => fifo_0_22_port, Y => data_out(22));
   U193 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_21_port, B1 => 
                           n43, B2 => fifo_0_21_port, Y => data_out(21));
   U194 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_20_port, B1 => 
                           n43, B2 => fifo_0_20_port, Y => data_out(20));
   U195 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_1_port, B1 => 
                           n43, B2 => fifo_0_1_port, Y => data_out(1));
   U196 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_19_port, B1 => 
                           n43, B2 => fifo_0_19_port, Y => data_out(19));
   U197 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_18_port, B1 => 
                           n43, B2 => fifo_0_18_port, Y => data_out(18));
   U198 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_17_port, B1 => 
                           n43, B2 => fifo_0_17_port, Y => data_out(17));
   U199 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_16_port, B1 => 
                           n43, B2 => fifo_0_16_port, Y => data_out(16));
   U200 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_15_port, B1 => 
                           n43, B2 => fifo_0_15_port, Y => data_out(15));
   U201 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_14_port, B1 => 
                           n43, B2 => fifo_0_14_port, Y => data_out(14));
   U202 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_13_port, B1 => 
                           n43, B2 => fifo_0_13_port, Y => data_out(13));
   U203 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_12_port, B1 => 
                           n43, B2 => fifo_0_12_port, Y => data_out(12));
   U204 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_11_port, B1 => 
                           n43, B2 => fifo_0_11_port, Y => data_out(11));
   U205 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_10_port, B1 => 
                           n43, B2 => fifo_0_10_port, Y => data_out(10));
   U206 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_0_port, B1 => 
                           n43, B2 => fifo_0_0_port, Y => data_out(0));
   U3 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n47, A2 => n238, B => 
                           valid_data_port, C => write_en, Y => n235);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_0_port, A2 => n17, B1 => 
                           data_in(0), B2 => n29, Y => n234);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_1_port, A2 => n17, B1 => 
                           data_in(1), B2 => n29, Y => n233);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_2_port, A2 => n17, B1 => 
                           data_in(2), B2 => n29, Y => n232);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_3_port, A2 => n17, B1 => 
                           data_in(3), B2 => n29, Y => n231);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_4_port, A2 => n17, B1 => 
                           data_in(4), B2 => n27, Y => n230);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_5_port, A2 => n17, B1 => 
                           data_in(5), B2 => n27, Y => n229);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_6_port, A2 => n17, B1 => 
                           data_in(6), B2 => n27, Y => n228);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_7_port, A2 => n17, B1 => 
                           data_in(7), B2 => n27, Y => n227);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_8_port, A2 => n17, B1 => 
                           data_in(8), B2 => n27, Y => n226);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_9_port, A2 => n17, B1 => 
                           data_in(9), B2 => n27, Y => n225);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_10_port, A2 => n17, B1 => 
                           data_in(10), B2 => n27, Y => n224);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_11_port, A2 => n17, B1 => 
                           data_in(11), B2 => n27, Y => n223);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_12_port, A2 => n17, B1 => 
                           data_in(12), B2 => n27, Y => n222);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_13_port, A2 => n17, B1 => 
                           data_in(13), B2 => n27, Y => n221);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_14_port, A2 => n17, B1 => 
                           data_in(14), B2 => n27, Y => n220);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_15_port, A2 => n17, B1 => 
                           data_in(15), B2 => n27, Y => n219);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_16_port, A2 => n17, B1 => 
                           data_in(16), B2 => n25, Y => n218);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_17_port, A2 => n17, B1 => 
                           data_in(17), B2 => n25, Y => n217);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_18_port, A2 => n17, B1 => 
                           data_in(18), B2 => n25, Y => n216);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_19_port, A2 => n17, B1 => 
                           data_in(19), B2 => n25, Y => n215);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_20_port, A2 => n17, B1 => 
                           data_in(20), B2 => n25, Y => n214);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_21_port, A2 => n17, B1 => 
                           data_in(21), B2 => n25, Y => n213);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_22_port, A2 => n17, B1 => 
                           data_in(22), B2 => n25, Y => n212);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_23_port, A2 => n17, B1 => 
                           data_in(23), B2 => n25, Y => n211);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_24_port, A2 => n17, B1 => 
                           data_in(24), B2 => n25, Y => n210);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_25_port, A2 => n17, B1 => 
                           data_in(25), B2 => n25, Y => n209);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_26_port, A2 => n17, B1 => 
                           data_in(26), B2 => n25, Y => n208);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_27_port, A2 => n17, B1 => 
                           data_in(27), B2 => n25, Y => n207);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_28_port, A2 => n17, B1 => 
                           data_in(28), B2 => n23, Y => n206);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_29_port, A2 => n17, B1 => 
                           data_in(29), B2 => n23, Y => n205);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_30_port, A2 => n17, B1 => 
                           data_in(30), B2 => n23, Y => n204);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_31_port, A2 => n17, B1 => 
                           data_in(31), B2 => n23, Y => n203);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_32_port, A2 => n17, B1 => 
                           data_in(32), B2 => n23, Y => n202);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_33_port, A2 => n17, B1 => 
                           data_in(33), B2 => n23, Y => n201);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_34_port, A2 => n17, B1 => 
                           data_in(34), B2 => n23, Y => n200);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_35_port, A2 => n17, B1 => 
                           data_in(35), B2 => n23, Y => n199);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_36_port, A2 => n17, B1 => 
                           data_in(36), B2 => n23, Y => n198);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_37_port, A2 => n17, B1 => 
                           data_in(37), B2 => n23, Y => n197);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_38_port, A2 => n17, B1 => 
                           data_in(38), B2 => n23, Y => n196);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_39_port, A2 => n17, B1 => 
                           data_in(39), B2 => n23, Y => n195);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_40_port, A2 => n17, B1 => 
                           data_in(40), B2 => n21, Y => n194);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_41_port, A2 => n17, B1 => 
                           data_in(41), B2 => n21, Y => n193);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_42_port, A2 => n17, B1 => 
                           data_in(42), B2 => n21, Y => n192);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_43_port, A2 => n17, B1 => 
                           data_in(43), B2 => n21, Y => n191);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_44_port, A2 => n17, B1 => 
                           data_in(44), B2 => n21, Y => n190);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_45_port, A2 => n17, B1 => 
                           data_in(45), B2 => n21, Y => n189);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_46_port, A2 => n17, B1 => 
                           data_in(46), B2 => n21, Y => n188);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_47_port, A2 => n17, B1 => 
                           data_in(47), B2 => n21, Y => n187);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_48_port, A2 => n17, B1 => 
                           data_in(48), B2 => n21, Y => n186);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_49_port, A2 => n17, B1 => 
                           data_in(49), B2 => n21, Y => n185);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_50_port, A2 => n17, B1 => 
                           data_in(50), B2 => n21, Y => n184);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_51_port, A2 => n17, B1 => 
                           data_in(51), B2 => n21, Y => n183);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_52_port, A2 => n17, B1 => 
                           data_in(52), B2 => n19, Y => n182);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_53_port, A2 => n17, B1 => 
                           data_in(53), B2 => n19, Y => n181);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_54_port, A2 => n17, B1 => 
                           data_in(54), B2 => n19, Y => n180);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_55_port, A2 => n17, B1 => 
                           data_in(55), B2 => n19, Y => n179);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_56_port, A2 => n17, B1 => 
                           data_in(56), B2 => n19, Y => n178);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_57_port, A2 => n17, B1 => 
                           data_in(57), B2 => n19, Y => n177);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_58_port, A2 => n17, B1 => 
                           data_in(58), B2 => n19, Y => n176);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_59_port, A2 => n17, B1 => 
                           data_in(59), B2 => n19, Y => n175);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_60_port, A2 => n17, B1 => 
                           data_in(60), B2 => n19, Y => n174);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_61_port, A2 => n17, B1 => 
                           data_in(61), B2 => n19, Y => n173);
   U67 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_62_port, A2 => n17, B1 => 
                           data_in(62), B2 => n19, Y => n172);
   U68 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_63_port, A2 => n17, B1 => 
                           data_in(63), B2 => n19, Y => n171);
   U70 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N9, Y => n237);
   U71 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_0_port, A2 => n3, B1 => 
                           data_in(0), B2 => n15, Y => n170);
   U72 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_1_port, A2 => n3, B1 => 
                           data_in(1), B2 => n15, Y => n169);
   U73 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_2_port, A2 => n3, B1 => 
                           data_in(2), B2 => n15, Y => n168);
   U74 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_3_port, A2 => n3, B1 => 
                           data_in(3), B2 => n15, Y => n167);
   U75 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_4_port, A2 => n3, B1 => 
                           data_in(4), B2 => n13, Y => n166);
   U76 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_5_port, A2 => n3, B1 => 
                           data_in(5), B2 => n13, Y => n165);
   U77 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_6_port, A2 => n3, B1 => 
                           data_in(6), B2 => n13, Y => n164);
   U78 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_7_port, A2 => n3, B1 => 
                           data_in(7), B2 => n13, Y => n163);
   U79 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_8_port, A2 => n3, B1 => 
                           data_in(8), B2 => n13, Y => n162);
   U80 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_9_port, A2 => n3, B1 => 
                           data_in(9), B2 => n13, Y => n161);
   U81 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_10_port, A2 => n3, B1 => 
                           data_in(10), B2 => n13, Y => n160);
   U82 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_11_port, A2 => n3, B1 => 
                           data_in(11), B2 => n13, Y => n159);
   U83 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_12_port, A2 => n3, B1 => 
                           data_in(12), B2 => n13, Y => n157);
   U84 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_13_port, A2 => n3, B1 => 
                           data_in(13), B2 => n13, Y => n155);
   U85 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_14_port, A2 => n3, B1 => 
                           data_in(14), B2 => n13, Y => n153);
   U86 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_15_port, A2 => n3, B1 => 
                           data_in(15), B2 => n13, Y => n151);
   U87 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_16_port, A2 => n3, B1 => 
                           data_in(16), B2 => n11, Y => n149);
   U88 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_17_port, A2 => n3, B1 => 
                           data_in(17), B2 => n11, Y => n147);
   U89 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_18_port, A2 => n3, B1 => 
                           data_in(18), B2 => n11, Y => n145);
   U90 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_19_port, A2 => n3, B1 => 
                           data_in(19), B2 => n11, Y => n143);
   U91 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_20_port, A2 => n3, B1 => 
                           data_in(20), B2 => n11, Y => n141);
   U92 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_21_port, A2 => n3, B1 => 
                           data_in(21), B2 => n11, Y => n139);
   U93 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_22_port, A2 => n3, B1 => 
                           data_in(22), B2 => n11, Y => n137);
   U94 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_23_port, A2 => n3, B1 => 
                           data_in(23), B2 => n11, Y => n135);
   U95 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_24_port, A2 => n3, B1 => 
                           data_in(24), B2 => n11, Y => n133);
   U96 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_25_port, A2 => n3, B1 => 
                           data_in(25), B2 => n11, Y => n131);
   U97 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_26_port, A2 => n3, B1 => 
                           data_in(26), B2 => n11, Y => n129);
   U98 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_27_port, A2 => n3, B1 => 
                           data_in(27), B2 => n11, Y => n127);
   U99 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_28_port, A2 => n3, B1 => 
                           data_in(28), B2 => n9_port, Y => n125);
   U100 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_29_port, A2 => n3, B1 => 
                           data_in(29), B2 => n9_port, Y => n123);
   U101 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_30_port, A2 => n3, B1 => 
                           data_in(30), B2 => n9_port, Y => n121);
   U102 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_31_port, A2 => n3, B1 => 
                           data_in(31), B2 => n9_port, Y => n119);
   U103 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_32_port, A2 => n3, B1 => 
                           data_in(32), B2 => n9_port, Y => n117);
   U104 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_33_port, A2 => n3, B1 => 
                           data_in(33), B2 => n9_port, Y => n115);
   U105 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_34_port, A2 => n3, B1 => 
                           data_in(34), B2 => n9_port, Y => n113);
   U106 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_35_port, A2 => n3, B1 => 
                           data_in(35), B2 => n9_port, Y => n111);
   U107 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_36_port, A2 => n3, B1 => 
                           data_in(36), B2 => n9_port, Y => n109);
   U108 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_37_port, A2 => n3, B1 => 
                           data_in(37), B2 => n9_port, Y => n107);
   U109 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_38_port, A2 => n3, B1 => 
                           data_in(38), B2 => n9_port, Y => n105);
   U110 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_39_port, A2 => n3, B1 => 
                           data_in(39), B2 => n9_port, Y => n103);
   U111 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_40_port, A2 => n3, B1 => 
                           data_in(40), B2 => n7_port, Y => n101);
   U112 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_41_port, A2 => n3, B1 => 
                           data_in(41), B2 => n7_port, Y => n99);
   U113 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_42_port, A2 => n3, B1 => 
                           data_in(42), B2 => n7_port, Y => n97);
   U114 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_43_port, A2 => n3, B1 => 
                           data_in(43), B2 => n7_port, Y => n95);
   U115 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_44_port, A2 => n3, B1 => 
                           data_in(44), B2 => n7_port, Y => n93);
   U116 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_45_port, A2 => n3, B1 => 
                           data_in(45), B2 => n7_port, Y => n91);
   U117 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_46_port, A2 => n3, B1 => 
                           data_in(46), B2 => n7_port, Y => n89);
   U118 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_47_port, A2 => n3, B1 => 
                           data_in(47), B2 => n7_port, Y => n87);
   U119 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_48_port, A2 => n3, B1 => 
                           data_in(48), B2 => n7_port, Y => n85);
   U120 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_49_port, A2 => n3, B1 => 
                           data_in(49), B2 => n7_port, Y => n83);
   U121 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_50_port, A2 => n3, B1 => 
                           data_in(50), B2 => n7_port, Y => n81);
   U122 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_51_port, A2 => n3, B1 => 
                           data_in(51), B2 => n7_port, Y => n79);
   U123 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_52_port, A2 => n3, B1 => 
                           data_in(52), B2 => n5, Y => n77);
   U124 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_53_port, A2 => n3, B1 => 
                           data_in(53), B2 => n5, Y => n75);
   U125 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_54_port, A2 => n3, B1 => 
                           data_in(54), B2 => n5, Y => n73);
   U126 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_55_port, A2 => n3, B1 => 
                           data_in(55), B2 => n5, Y => n71);
   U127 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_56_port, A2 => n3, B1 => 
                           data_in(56), B2 => n5, Y => n69);
   U128 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_57_port, A2 => n3, B1 => 
                           data_in(57), B2 => n5, Y => n67);
   U129 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_58_port, A2 => n3, B1 => 
                           data_in(58), B2 => n5, Y => n65);
   U130 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_59_port, A2 => n3, B1 => 
                           data_in(59), B2 => n5, Y => n63);
   U131 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_60_port, A2 => n3, B1 => 
                           data_in(60), B2 => n5, Y => n61);
   U132 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_61_port, A2 => n3, B1 => 
                           data_in(61), B2 => n5, Y => n59);
   U133 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_62_port, A2 => n3, B1 => 
                           data_in(62), B2 => n5, Y => n57);
   U134 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_63_port, A2 => n3, B1 => 
                           data_in(63), B2 => n5, Y => n55);
   U136 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N7, Y => n236);
   U137 : OAI22xp5_ASAP7_75t_R port map( A1 => n31, A2 => read_en, B1 => n43, 
                           B2 => n47, Y => n53);
   U139 : OAI22xp5_ASAP7_75t_R port map( A1 => N9, A2 => n49, B1 => write_en, 
                           B2 => N7, Y => n51);
   write_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK 
                           => clk, RESET => n45, SET => n1, QN => N7);
   fifo_reg_1_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n55, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_63_port);
   fifo_reg_1_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n57, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_62_port);
   fifo_reg_1_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n59, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_61_port);
   fifo_reg_1_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n61, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_60_port);
   fifo_reg_0_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n171, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_63_port);
   fifo_reg_0_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n172, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_62_port);
   fifo_reg_0_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n173, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_61_port);
   fifo_reg_0_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n174, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_60_port);
   fifo_reg_1_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n167, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_3_port);
   fifo_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n168, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_2_port);
   fifo_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n169, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_1_port);
   fifo_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n170, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_0_port);
   fifo_reg_1_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n63, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_59_port);
   fifo_reg_1_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n65, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_58_port);
   fifo_reg_1_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n67, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_57_port);
   fifo_reg_1_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n69, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_56_port);
   fifo_reg_1_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n71, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_55_port);
   fifo_reg_1_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n73, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_54_port);
   fifo_reg_1_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n75, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_53_port);
   fifo_reg_1_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n77, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_52_port);
   fifo_reg_1_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_51_port);
   fifo_reg_1_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_50_port);
   fifo_reg_1_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_49_port);
   fifo_reg_1_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_48_port);
   fifo_reg_1_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_47_port);
   fifo_reg_1_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_46_port);
   fifo_reg_1_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_45_port);
   fifo_reg_1_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_44_port);
   fifo_reg_1_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_43_port);
   fifo_reg_1_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_42_port);
   fifo_reg_1_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_41_port);
   fifo_reg_1_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_40_port);
   fifo_reg_1_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_39_port);
   fifo_reg_1_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_38_port);
   fifo_reg_1_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_37_port);
   fifo_reg_1_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_36_port);
   fifo_reg_1_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_35_port);
   fifo_reg_1_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_34_port);
   fifo_reg_1_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n115, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_33_port);
   fifo_reg_1_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n117, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_32_port);
   fifo_reg_1_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n119, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_31_port);
   fifo_reg_1_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n121, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_30_port);
   fifo_reg_1_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n123, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_29_port);
   fifo_reg_1_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n125, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_28_port);
   fifo_reg_1_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n127, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_27_port);
   fifo_reg_1_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n129, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_26_port);
   fifo_reg_1_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n131, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_25_port);
   fifo_reg_1_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n133, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_24_port);
   fifo_reg_1_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n135, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_23_port);
   fifo_reg_1_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n137, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_22_port);
   fifo_reg_1_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n139, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_21_port);
   fifo_reg_1_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n141, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_20_port);
   fifo_reg_1_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n143, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_19_port);
   fifo_reg_1_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n145, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_18_port);
   fifo_reg_1_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n147, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_17_port);
   fifo_reg_1_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n149, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_16_port);
   fifo_reg_1_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n151, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_15_port);
   fifo_reg_1_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n153, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_14_port);
   fifo_reg_1_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n155, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_13_port);
   fifo_reg_1_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n157, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_12_port);
   fifo_reg_1_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n159, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_11_port);
   fifo_reg_1_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n160, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_10_port);
   fifo_reg_1_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n161, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_9_port);
   fifo_reg_1_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n162, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_8_port);
   fifo_reg_1_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n163, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_7_port);
   fifo_reg_1_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n164, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_6_port);
   fifo_reg_1_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n165, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_5_port);
   fifo_reg_1_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n166, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_4_port);
   fifo_reg_0_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n231, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_3_port);
   fifo_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n232, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_2_port);
   fifo_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n233, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_1_port);
   fifo_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n234, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_0_port);
   fifo_reg_0_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n175, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_59_port);
   fifo_reg_0_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n176, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_58_port);
   fifo_reg_0_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n177, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_57_port);
   fifo_reg_0_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n178, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_56_port);
   fifo_reg_0_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n179, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_55_port);
   fifo_reg_0_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n180, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_54_port);
   fifo_reg_0_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n181, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_53_port);
   fifo_reg_0_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n182, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_52_port);
   fifo_reg_0_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n183, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_51_port);
   fifo_reg_0_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n184, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_50_port);
   fifo_reg_0_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n185, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_49_port);
   fifo_reg_0_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n186, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_48_port);
   fifo_reg_0_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n187, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_47_port);
   fifo_reg_0_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n188, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_46_port);
   fifo_reg_0_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n189, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_45_port);
   fifo_reg_0_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n190, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_44_port);
   fifo_reg_0_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n191, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_43_port);
   fifo_reg_0_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n192, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_42_port);
   fifo_reg_0_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n193, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_41_port);
   fifo_reg_0_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n194, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_40_port);
   fifo_reg_0_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n195, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_39_port);
   fifo_reg_0_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n196, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_38_port);
   fifo_reg_0_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n197, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_37_port);
   fifo_reg_0_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n198, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_36_port);
   fifo_reg_0_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n199, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_35_port);
   fifo_reg_0_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n200, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_34_port);
   fifo_reg_0_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n201, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_33_port);
   fifo_reg_0_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n202, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_32_port);
   fifo_reg_0_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n203, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_31_port);
   fifo_reg_0_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n204, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_30_port);
   fifo_reg_0_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n205, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_29_port);
   fifo_reg_0_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n206, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_28_port);
   fifo_reg_0_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n207, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_27_port);
   fifo_reg_0_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n208, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_26_port);
   fifo_reg_0_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n209, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_25_port);
   fifo_reg_0_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n210, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_24_port);
   fifo_reg_0_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n211, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_23_port);
   fifo_reg_0_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n212, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_22_port);
   fifo_reg_0_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n213, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_21_port);
   fifo_reg_0_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n214, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_20_port);
   fifo_reg_0_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n215, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_19_port);
   fifo_reg_0_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n216, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_18_port);
   fifo_reg_0_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n217, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_17_port);
   fifo_reg_0_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n218, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_16_port);
   fifo_reg_0_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n219, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_15_port);
   fifo_reg_0_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n220, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_14_port);
   fifo_reg_0_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n221, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_13_port);
   fifo_reg_0_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n222, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_12_port);
   fifo_reg_0_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n223, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_11_port);
   fifo_reg_0_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n224, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_10_port);
   fifo_reg_0_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n225, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_9_port);
   fifo_reg_0_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n226, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_8_port);
   fifo_reg_0_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n227, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_7_port);
   fifo_reg_0_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n228, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_6_port);
   fifo_reg_0_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n229, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_5_port);
   fifo_reg_0_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n230, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_4_port);
   read_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK 
                           => clk, RESET => n45, SET => n1, QN => 
                           read_pointer_0_port);
   valid_data_reg : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n235, CLK => clk, 
                           RESET => n45, SET => n1, QN => valid_data_port);
   U69 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U135 : INVx3_ASAP7_75t_R port map( A => rst, Y => n45);
   U138 : INVx1_ASAP7_75t_R port map( A => n29, Y => n17);
   U140 : INVx1_ASAP7_75t_R port map( A => n15, Y => n3);
   U141 : INVx1_ASAP7_75t_R port map( A => n31, Y => n43);
   U142 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n29);
   U207 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n15);
   U208 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n27);
   U209 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n25);
   U210 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n23);
   U211 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n21);
   U212 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n19);
   U213 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n13);
   U214 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n11);
   U215 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n9_port);
   U216 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n7_port);
   U217 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n5);
   U218 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n31);
   U219 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n33);
   U220 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n41);
   U221 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n39);
   U222 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n37);
   U223 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n35);
   U224 : INVx1_ASAP7_75t_R port map( A => read_en, Y => n47);
   U225 : INVx1_ASAP7_75t_R port map( A => N7, Y => N9);
   U226 : INVx1_ASAP7_75t_R port map( A => write_en, Y => n49);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity fifo_buff_depth2_11 is

   port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, clk, 
         rst : in std_logic;  data_out : out std_logic_vector (63 downto 0);  
         valid_data : out std_logic);

end fifo_buff_depth2_11;

architecture SYN_rtl of fifo_buff_depth2_11 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx3_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal valid_data_port, read_pointer_0_port, fifo_1_63_port, fifo_1_62_port,
      fifo_1_61_port, fifo_1_60_port, fifo_1_59_port, fifo_1_58_port, 
      fifo_1_57_port, fifo_1_56_port, fifo_1_55_port, fifo_1_54_port, 
      fifo_1_53_port, fifo_1_52_port, fifo_1_51_port, fifo_1_50_port, 
      fifo_1_49_port, fifo_1_48_port, fifo_1_47_port, fifo_1_46_port, 
      fifo_1_45_port, fifo_1_44_port, fifo_1_43_port, fifo_1_42_port, 
      fifo_1_41_port, fifo_1_40_port, fifo_1_39_port, fifo_1_38_port, 
      fifo_1_37_port, fifo_1_36_port, fifo_1_35_port, fifo_1_34_port, 
      fifo_1_33_port, fifo_1_32_port, fifo_1_31_port, fifo_1_30_port, 
      fifo_1_29_port, fifo_1_28_port, fifo_1_27_port, fifo_1_26_port, 
      fifo_1_25_port, fifo_1_24_port, fifo_1_23_port, fifo_1_22_port, 
      fifo_1_21_port, fifo_1_20_port, fifo_1_19_port, fifo_1_18_port, 
      fifo_1_17_port, fifo_1_16_port, fifo_1_15_port, fifo_1_14_port, 
      fifo_1_13_port, fifo_1_12_port, fifo_1_11_port, fifo_1_10_port, 
      fifo_1_9_port, fifo_1_8_port, fifo_1_7_port, fifo_1_6_port, fifo_1_5_port
      , fifo_1_4_port, fifo_1_3_port, fifo_1_2_port, fifo_1_1_port, 
      fifo_1_0_port, fifo_0_63_port, fifo_0_62_port, fifo_0_61_port, 
      fifo_0_60_port, fifo_0_59_port, fifo_0_58_port, fifo_0_57_port, 
      fifo_0_56_port, fifo_0_55_port, fifo_0_54_port, fifo_0_53_port, 
      fifo_0_52_port, fifo_0_51_port, fifo_0_50_port, fifo_0_49_port, 
      fifo_0_48_port, fifo_0_47_port, fifo_0_46_port, fifo_0_45_port, 
      fifo_0_44_port, fifo_0_43_port, fifo_0_42_port, fifo_0_41_port, 
      fifo_0_40_port, fifo_0_39_port, fifo_0_38_port, fifo_0_37_port, 
      fifo_0_36_port, fifo_0_35_port, fifo_0_34_port, fifo_0_33_port, 
      fifo_0_32_port, fifo_0_31_port, fifo_0_30_port, fifo_0_29_port, 
      fifo_0_28_port, fifo_0_27_port, fifo_0_26_port, fifo_0_25_port, 
      fifo_0_24_port, fifo_0_23_port, fifo_0_22_port, fifo_0_21_port, 
      fifo_0_20_port, fifo_0_19_port, fifo_0_18_port, fifo_0_17_port, 
      fifo_0_16_port, fifo_0_15_port, fifo_0_14_port, fifo_0_13_port, 
      fifo_0_12_port, fifo_0_11_port, fifo_0_10_port, fifo_0_9_port, 
      fifo_0_8_port, fifo_0_7_port, fifo_0_6_port, fifo_0_5_port, fifo_0_4_port
      , fifo_0_3_port, fifo_0_2_port, fifo_0_1_port, fifo_0_0_port, N7, N9, n1,
      n3, n5, n7_port, n9_port, n11, n13, n15, n17, n19, n21, n23, n25, n27, 
      n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57
      , n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, 
      n87, n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, n111, 
      n113, n115, n117, n119, n121, n123, n125, n127, n129, n131, n133, n135, 
      n137, n139, n141, n143, n145, n147, n149, n151, n153, n155, n157, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238 : std_logic;

begin
   valid_data <= valid_data_port;
   
   U4 : XOR2xp5_ASAP7_75t_R port map( A => N7, B => n43, Y => n238);
   U143 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_9_port, B1 => 
                           n43, B2 => fifo_0_9_port, Y => data_out(9));
   U144 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_8_port, B1 => 
                           n43, B2 => fifo_0_8_port, Y => data_out(8));
   U145 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_7_port, B1 => 
                           n43, B2 => fifo_0_7_port, Y => data_out(7));
   U146 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_6_port, B1 => 
                           n43, B2 => fifo_0_6_port, Y => data_out(6));
   U147 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_63_port, B1 => 
                           n43, B2 => fifo_0_63_port, Y => data_out(63));
   U148 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_62_port, B1 => 
                           n43, B2 => fifo_0_62_port, Y => data_out(62));
   U149 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_61_port, B1 => 
                           n43, B2 => fifo_0_61_port, Y => data_out(61));
   U150 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_60_port, B1 => 
                           n43, B2 => fifo_0_60_port, Y => data_out(60));
   U151 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_5_port, B1 => 
                           n43, B2 => fifo_0_5_port, Y => data_out(5));
   U152 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_59_port, B1 => 
                           n43, B2 => fifo_0_59_port, Y => data_out(59));
   U153 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_58_port, B1 => 
                           n43, B2 => fifo_0_58_port, Y => data_out(58));
   U154 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_57_port, B1 => 
                           n43, B2 => fifo_0_57_port, Y => data_out(57));
   U155 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_56_port, B1 => 
                           n43, B2 => fifo_0_56_port, Y => data_out(56));
   U156 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_55_port, B1 => 
                           n43, B2 => fifo_0_55_port, Y => data_out(55));
   U157 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_54_port, B1 => 
                           n43, B2 => fifo_0_54_port, Y => data_out(54));
   U158 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_53_port, B1 => 
                           n43, B2 => fifo_0_53_port, Y => data_out(53));
   U159 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_52_port, B1 => 
                           n43, B2 => fifo_0_52_port, Y => data_out(52));
   U160 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_51_port, B1 => 
                           n43, B2 => fifo_0_51_port, Y => data_out(51));
   U161 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_50_port, B1 => 
                           n43, B2 => fifo_0_50_port, Y => data_out(50));
   U162 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_4_port, B1 => 
                           n43, B2 => fifo_0_4_port, Y => data_out(4));
   U163 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_49_port, B1 => 
                           n43, B2 => fifo_0_49_port, Y => data_out(49));
   U164 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_48_port, B1 => 
                           n43, B2 => fifo_0_48_port, Y => data_out(48));
   U165 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_47_port, B1 => 
                           n43, B2 => fifo_0_47_port, Y => data_out(47));
   U166 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_46_port, B1 => 
                           n43, B2 => fifo_0_46_port, Y => data_out(46));
   U167 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_45_port, B1 => 
                           n43, B2 => fifo_0_45_port, Y => data_out(45));
   U168 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_44_port, B1 => 
                           n43, B2 => fifo_0_44_port, Y => data_out(44));
   U169 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_43_port, B1 => 
                           n43, B2 => fifo_0_43_port, Y => data_out(43));
   U170 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_42_port, B1 => 
                           n43, B2 => fifo_0_42_port, Y => data_out(42));
   U171 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_41_port, B1 => 
                           n43, B2 => fifo_0_41_port, Y => data_out(41));
   U172 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_40_port, B1 => 
                           n43, B2 => fifo_0_40_port, Y => data_out(40));
   U173 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_3_port, B1 => 
                           n43, B2 => fifo_0_3_port, Y => data_out(3));
   U174 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_39_port, B1 => 
                           n43, B2 => fifo_0_39_port, Y => data_out(39));
   U175 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_38_port, B1 => 
                           n43, B2 => fifo_0_38_port, Y => data_out(38));
   U176 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_37_port, B1 => 
                           n43, B2 => fifo_0_37_port, Y => data_out(37));
   U177 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_36_port, B1 => 
                           n43, B2 => fifo_0_36_port, Y => data_out(36));
   U178 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_35_port, B1 => 
                           n43, B2 => fifo_0_35_port, Y => data_out(35));
   U179 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_34_port, B1 => 
                           n43, B2 => fifo_0_34_port, Y => data_out(34));
   U180 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_33_port, B1 => 
                           n43, B2 => fifo_0_33_port, Y => data_out(33));
   U181 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_32_port, B1 => 
                           n43, B2 => fifo_0_32_port, Y => data_out(32));
   U182 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_31_port, B1 => 
                           n43, B2 => fifo_0_31_port, Y => data_out(31));
   U183 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_30_port, B1 => 
                           n43, B2 => fifo_0_30_port, Y => data_out(30));
   U184 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_2_port, B1 => 
                           n43, B2 => fifo_0_2_port, Y => data_out(2));
   U185 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_29_port, B1 => 
                           n43, B2 => fifo_0_29_port, Y => data_out(29));
   U186 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_28_port, B1 => 
                           n43, B2 => fifo_0_28_port, Y => data_out(28));
   U187 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_27_port, B1 => 
                           n43, B2 => fifo_0_27_port, Y => data_out(27));
   U188 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_26_port, B1 => 
                           n43, B2 => fifo_0_26_port, Y => data_out(26));
   U189 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_25_port, B1 => 
                           n43, B2 => fifo_0_25_port, Y => data_out(25));
   U190 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_24_port, B1 => 
                           n43, B2 => fifo_0_24_port, Y => data_out(24));
   U191 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_23_port, B1 => 
                           n43, B2 => fifo_0_23_port, Y => data_out(23));
   U192 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_22_port, B1 => 
                           n43, B2 => fifo_0_22_port, Y => data_out(22));
   U193 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_21_port, B1 => 
                           n43, B2 => fifo_0_21_port, Y => data_out(21));
   U194 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_20_port, B1 => 
                           n43, B2 => fifo_0_20_port, Y => data_out(20));
   U195 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_1_port, B1 => 
                           n43, B2 => fifo_0_1_port, Y => data_out(1));
   U196 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_19_port, B1 => 
                           n43, B2 => fifo_0_19_port, Y => data_out(19));
   U197 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_18_port, B1 => 
                           n43, B2 => fifo_0_18_port, Y => data_out(18));
   U198 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_17_port, B1 => 
                           n43, B2 => fifo_0_17_port, Y => data_out(17));
   U199 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_16_port, B1 => 
                           n43, B2 => fifo_0_16_port, Y => data_out(16));
   U200 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_15_port, B1 => 
                           n43, B2 => fifo_0_15_port, Y => data_out(15));
   U201 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_14_port, B1 => 
                           n43, B2 => fifo_0_14_port, Y => data_out(14));
   U202 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_13_port, B1 => 
                           n43, B2 => fifo_0_13_port, Y => data_out(13));
   U203 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_12_port, B1 => 
                           n43, B2 => fifo_0_12_port, Y => data_out(12));
   U204 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_11_port, B1 => 
                           n43, B2 => fifo_0_11_port, Y => data_out(11));
   U205 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_10_port, B1 => 
                           n43, B2 => fifo_0_10_port, Y => data_out(10));
   U206 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_0_port, B1 => 
                           n43, B2 => fifo_0_0_port, Y => data_out(0));
   U3 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n45, A2 => n238, B => 
                           valid_data_port, C => write_en, Y => n235);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_0_port, A2 => n17, B1 => 
                           data_in(0), B2 => n29, Y => n234);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_1_port, A2 => n17, B1 => 
                           data_in(1), B2 => n29, Y => n233);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_2_port, A2 => n17, B1 => 
                           data_in(2), B2 => n29, Y => n232);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_3_port, A2 => n17, B1 => 
                           data_in(3), B2 => n29, Y => n231);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_4_port, A2 => n17, B1 => 
                           data_in(4), B2 => n27, Y => n230);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_5_port, A2 => n17, B1 => 
                           data_in(5), B2 => n27, Y => n229);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_6_port, A2 => n17, B1 => 
                           data_in(6), B2 => n27, Y => n228);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_7_port, A2 => n17, B1 => 
                           data_in(7), B2 => n27, Y => n227);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_8_port, A2 => n17, B1 => 
                           data_in(8), B2 => n27, Y => n226);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_9_port, A2 => n17, B1 => 
                           data_in(9), B2 => n27, Y => n225);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_10_port, A2 => n17, B1 => 
                           data_in(10), B2 => n27, Y => n224);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_11_port, A2 => n17, B1 => 
                           data_in(11), B2 => n27, Y => n223);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_12_port, A2 => n17, B1 => 
                           data_in(12), B2 => n27, Y => n222);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_13_port, A2 => n17, B1 => 
                           data_in(13), B2 => n27, Y => n221);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_14_port, A2 => n17, B1 => 
                           data_in(14), B2 => n27, Y => n220);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_15_port, A2 => n17, B1 => 
                           data_in(15), B2 => n27, Y => n219);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_16_port, A2 => n17, B1 => 
                           data_in(16), B2 => n25, Y => n218);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_17_port, A2 => n17, B1 => 
                           data_in(17), B2 => n25, Y => n217);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_18_port, A2 => n17, B1 => 
                           data_in(18), B2 => n25, Y => n216);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_19_port, A2 => n17, B1 => 
                           data_in(19), B2 => n25, Y => n215);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_20_port, A2 => n17, B1 => 
                           data_in(20), B2 => n25, Y => n214);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_21_port, A2 => n17, B1 => 
                           data_in(21), B2 => n25, Y => n213);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_22_port, A2 => n17, B1 => 
                           data_in(22), B2 => n25, Y => n212);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_23_port, A2 => n17, B1 => 
                           data_in(23), B2 => n25, Y => n211);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_24_port, A2 => n17, B1 => 
                           data_in(24), B2 => n25, Y => n210);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_25_port, A2 => n17, B1 => 
                           data_in(25), B2 => n25, Y => n209);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_26_port, A2 => n17, B1 => 
                           data_in(26), B2 => n25, Y => n208);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_27_port, A2 => n17, B1 => 
                           data_in(27), B2 => n25, Y => n207);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_28_port, A2 => n17, B1 => 
                           data_in(28), B2 => n23, Y => n206);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_29_port, A2 => n17, B1 => 
                           data_in(29), B2 => n23, Y => n205);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_30_port, A2 => n17, B1 => 
                           data_in(30), B2 => n23, Y => n204);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_31_port, A2 => n17, B1 => 
                           data_in(31), B2 => n23, Y => n203);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_32_port, A2 => n17, B1 => 
                           data_in(32), B2 => n23, Y => n202);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_33_port, A2 => n17, B1 => 
                           data_in(33), B2 => n23, Y => n201);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_34_port, A2 => n17, B1 => 
                           data_in(34), B2 => n23, Y => n200);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_35_port, A2 => n17, B1 => 
                           data_in(35), B2 => n23, Y => n199);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_36_port, A2 => n17, B1 => 
                           data_in(36), B2 => n23, Y => n198);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_37_port, A2 => n17, B1 => 
                           data_in(37), B2 => n23, Y => n197);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_38_port, A2 => n17, B1 => 
                           data_in(38), B2 => n23, Y => n196);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_39_port, A2 => n17, B1 => 
                           data_in(39), B2 => n23, Y => n195);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_40_port, A2 => n17, B1 => 
                           data_in(40), B2 => n21, Y => n194);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_41_port, A2 => n17, B1 => 
                           data_in(41), B2 => n21, Y => n193);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_42_port, A2 => n17, B1 => 
                           data_in(42), B2 => n21, Y => n192);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_43_port, A2 => n17, B1 => 
                           data_in(43), B2 => n21, Y => n191);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_44_port, A2 => n17, B1 => 
                           data_in(44), B2 => n21, Y => n190);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_45_port, A2 => n17, B1 => 
                           data_in(45), B2 => n21, Y => n189);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_46_port, A2 => n17, B1 => 
                           data_in(46), B2 => n21, Y => n188);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_47_port, A2 => n17, B1 => 
                           data_in(47), B2 => n21, Y => n187);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_48_port, A2 => n17, B1 => 
                           data_in(48), B2 => n21, Y => n186);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_49_port, A2 => n17, B1 => 
                           data_in(49), B2 => n21, Y => n185);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_50_port, A2 => n17, B1 => 
                           data_in(50), B2 => n21, Y => n184);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_51_port, A2 => n17, B1 => 
                           data_in(51), B2 => n21, Y => n183);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_52_port, A2 => n17, B1 => 
                           data_in(52), B2 => n19, Y => n182);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_53_port, A2 => n17, B1 => 
                           data_in(53), B2 => n19, Y => n181);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_54_port, A2 => n17, B1 => 
                           data_in(54), B2 => n19, Y => n180);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_55_port, A2 => n17, B1 => 
                           data_in(55), B2 => n19, Y => n179);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_56_port, A2 => n17, B1 => 
                           data_in(56), B2 => n19, Y => n178);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_57_port, A2 => n17, B1 => 
                           data_in(57), B2 => n19, Y => n177);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_58_port, A2 => n17, B1 => 
                           data_in(58), B2 => n19, Y => n176);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_59_port, A2 => n17, B1 => 
                           data_in(59), B2 => n19, Y => n175);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_60_port, A2 => n17, B1 => 
                           data_in(60), B2 => n19, Y => n174);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_61_port, A2 => n17, B1 => 
                           data_in(61), B2 => n19, Y => n173);
   U67 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_62_port, A2 => n17, B1 => 
                           data_in(62), B2 => n19, Y => n172);
   U68 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_63_port, A2 => n17, B1 => 
                           data_in(63), B2 => n19, Y => n171);
   U70 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N9, Y => n237);
   U71 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_0_port, A2 => n3, B1 => 
                           data_in(0), B2 => n15, Y => n170);
   U72 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_1_port, A2 => n3, B1 => 
                           data_in(1), B2 => n15, Y => n169);
   U73 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_2_port, A2 => n3, B1 => 
                           data_in(2), B2 => n15, Y => n168);
   U74 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_3_port, A2 => n3, B1 => 
                           data_in(3), B2 => n15, Y => n167);
   U75 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_4_port, A2 => n3, B1 => 
                           data_in(4), B2 => n13, Y => n166);
   U76 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_5_port, A2 => n3, B1 => 
                           data_in(5), B2 => n13, Y => n165);
   U77 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_6_port, A2 => n3, B1 => 
                           data_in(6), B2 => n13, Y => n164);
   U78 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_7_port, A2 => n3, B1 => 
                           data_in(7), B2 => n13, Y => n163);
   U79 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_8_port, A2 => n3, B1 => 
                           data_in(8), B2 => n13, Y => n162);
   U80 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_9_port, A2 => n3, B1 => 
                           data_in(9), B2 => n13, Y => n161);
   U81 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_10_port, A2 => n3, B1 => 
                           data_in(10), B2 => n13, Y => n160);
   U82 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_11_port, A2 => n3, B1 => 
                           data_in(11), B2 => n13, Y => n159);
   U83 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_12_port, A2 => n3, B1 => 
                           data_in(12), B2 => n13, Y => n157);
   U84 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_13_port, A2 => n3, B1 => 
                           data_in(13), B2 => n13, Y => n155);
   U85 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_14_port, A2 => n3, B1 => 
                           data_in(14), B2 => n13, Y => n153);
   U86 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_15_port, A2 => n3, B1 => 
                           data_in(15), B2 => n13, Y => n151);
   U87 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_16_port, A2 => n3, B1 => 
                           data_in(16), B2 => n11, Y => n149);
   U88 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_17_port, A2 => n3, B1 => 
                           data_in(17), B2 => n11, Y => n147);
   U89 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_18_port, A2 => n3, B1 => 
                           data_in(18), B2 => n11, Y => n145);
   U90 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_19_port, A2 => n3, B1 => 
                           data_in(19), B2 => n11, Y => n143);
   U91 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_20_port, A2 => n3, B1 => 
                           data_in(20), B2 => n11, Y => n141);
   U92 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_21_port, A2 => n3, B1 => 
                           data_in(21), B2 => n11, Y => n139);
   U93 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_22_port, A2 => n3, B1 => 
                           data_in(22), B2 => n11, Y => n137);
   U94 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_23_port, A2 => n3, B1 => 
                           data_in(23), B2 => n11, Y => n135);
   U95 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_24_port, A2 => n3, B1 => 
                           data_in(24), B2 => n11, Y => n133);
   U96 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_25_port, A2 => n3, B1 => 
                           data_in(25), B2 => n11, Y => n131);
   U97 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_26_port, A2 => n3, B1 => 
                           data_in(26), B2 => n11, Y => n129);
   U98 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_27_port, A2 => n3, B1 => 
                           data_in(27), B2 => n11, Y => n127);
   U99 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_28_port, A2 => n3, B1 => 
                           data_in(28), B2 => n9_port, Y => n125);
   U100 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_29_port, A2 => n3, B1 => 
                           data_in(29), B2 => n9_port, Y => n123);
   U101 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_30_port, A2 => n3, B1 => 
                           data_in(30), B2 => n9_port, Y => n121);
   U102 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_31_port, A2 => n3, B1 => 
                           data_in(31), B2 => n9_port, Y => n119);
   U103 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_32_port, A2 => n3, B1 => 
                           data_in(32), B2 => n9_port, Y => n117);
   U104 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_33_port, A2 => n3, B1 => 
                           data_in(33), B2 => n9_port, Y => n115);
   U105 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_34_port, A2 => n3, B1 => 
                           data_in(34), B2 => n9_port, Y => n113);
   U106 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_35_port, A2 => n3, B1 => 
                           data_in(35), B2 => n9_port, Y => n111);
   U107 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_36_port, A2 => n3, B1 => 
                           data_in(36), B2 => n9_port, Y => n109);
   U108 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_37_port, A2 => n3, B1 => 
                           data_in(37), B2 => n9_port, Y => n107);
   U109 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_38_port, A2 => n3, B1 => 
                           data_in(38), B2 => n9_port, Y => n105);
   U110 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_39_port, A2 => n3, B1 => 
                           data_in(39), B2 => n9_port, Y => n103);
   U111 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_40_port, A2 => n3, B1 => 
                           data_in(40), B2 => n7_port, Y => n101);
   U112 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_41_port, A2 => n3, B1 => 
                           data_in(41), B2 => n7_port, Y => n99);
   U113 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_42_port, A2 => n3, B1 => 
                           data_in(42), B2 => n7_port, Y => n97);
   U114 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_43_port, A2 => n3, B1 => 
                           data_in(43), B2 => n7_port, Y => n95);
   U115 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_44_port, A2 => n3, B1 => 
                           data_in(44), B2 => n7_port, Y => n93);
   U116 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_45_port, A2 => n3, B1 => 
                           data_in(45), B2 => n7_port, Y => n91);
   U117 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_46_port, A2 => n3, B1 => 
                           data_in(46), B2 => n7_port, Y => n89);
   U118 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_47_port, A2 => n3, B1 => 
                           data_in(47), B2 => n7_port, Y => n87);
   U119 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_48_port, A2 => n3, B1 => 
                           data_in(48), B2 => n7_port, Y => n85);
   U120 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_49_port, A2 => n3, B1 => 
                           data_in(49), B2 => n7_port, Y => n83);
   U121 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_50_port, A2 => n3, B1 => 
                           data_in(50), B2 => n7_port, Y => n81);
   U122 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_51_port, A2 => n3, B1 => 
                           data_in(51), B2 => n7_port, Y => n79);
   U123 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_52_port, A2 => n3, B1 => 
                           data_in(52), B2 => n5, Y => n77);
   U124 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_53_port, A2 => n3, B1 => 
                           data_in(53), B2 => n5, Y => n75);
   U125 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_54_port, A2 => n3, B1 => 
                           data_in(54), B2 => n5, Y => n73);
   U126 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_55_port, A2 => n3, B1 => 
                           data_in(55), B2 => n5, Y => n71);
   U127 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_56_port, A2 => n3, B1 => 
                           data_in(56), B2 => n5, Y => n69);
   U128 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_57_port, A2 => n3, B1 => 
                           data_in(57), B2 => n5, Y => n67);
   U129 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_58_port, A2 => n3, B1 => 
                           data_in(58), B2 => n5, Y => n65);
   U130 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_59_port, A2 => n3, B1 => 
                           data_in(59), B2 => n5, Y => n63);
   U131 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_60_port, A2 => n3, B1 => 
                           data_in(60), B2 => n5, Y => n61);
   U132 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_61_port, A2 => n3, B1 => 
                           data_in(61), B2 => n5, Y => n59);
   U133 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_62_port, A2 => n3, B1 => 
                           data_in(62), B2 => n5, Y => n57);
   U134 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_63_port, A2 => n3, B1 => 
                           data_in(63), B2 => n5, Y => n55);
   U136 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N7, Y => n236);
   U137 : OAI22xp5_ASAP7_75t_R port map( A1 => n31, A2 => read_en, B1 => n43, 
                           B2 => n45, Y => n53);
   U139 : OAI22xp5_ASAP7_75t_R port map( A1 => N9, A2 => n49, B1 => write_en, 
                           B2 => N7, Y => n51);
   write_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK 
                           => clk, RESET => n47, SET => n1, QN => N7);
   fifo_reg_1_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n55, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_63_port);
   fifo_reg_1_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n57, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_62_port);
   fifo_reg_1_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n59, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_61_port);
   fifo_reg_1_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n61, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_60_port);
   fifo_reg_0_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n171, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_63_port);
   fifo_reg_0_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n172, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_62_port);
   fifo_reg_0_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n173, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_61_port);
   fifo_reg_0_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n174, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_60_port);
   fifo_reg_1_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n167, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_3_port);
   fifo_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n168, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_2_port);
   fifo_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n169, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_1_port);
   fifo_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n170, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_0_port);
   fifo_reg_1_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n63, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_59_port);
   fifo_reg_1_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n65, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_58_port);
   fifo_reg_1_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n67, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_57_port);
   fifo_reg_1_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n69, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_56_port);
   fifo_reg_1_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n71, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_55_port);
   fifo_reg_1_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n73, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_54_port);
   fifo_reg_1_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n75, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_53_port);
   fifo_reg_1_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n77, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_52_port);
   fifo_reg_1_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_51_port);
   fifo_reg_1_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_50_port);
   fifo_reg_1_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_49_port);
   fifo_reg_1_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_48_port);
   fifo_reg_1_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_47_port);
   fifo_reg_1_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_46_port);
   fifo_reg_1_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_45_port);
   fifo_reg_1_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_44_port);
   fifo_reg_1_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_43_port);
   fifo_reg_1_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_42_port);
   fifo_reg_1_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_41_port);
   fifo_reg_1_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_40_port);
   fifo_reg_1_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_39_port);
   fifo_reg_1_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_38_port);
   fifo_reg_1_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_37_port);
   fifo_reg_1_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_36_port);
   fifo_reg_1_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_35_port);
   fifo_reg_1_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_34_port);
   fifo_reg_1_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n115, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_33_port);
   fifo_reg_1_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n117, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_32_port);
   fifo_reg_1_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n119, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_31_port);
   fifo_reg_1_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n121, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_30_port);
   fifo_reg_1_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n123, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_29_port);
   fifo_reg_1_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n125, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_28_port);
   fifo_reg_1_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n127, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_27_port);
   fifo_reg_1_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n129, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_26_port);
   fifo_reg_1_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n131, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_25_port);
   fifo_reg_1_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n133, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_24_port);
   fifo_reg_1_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n135, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_23_port);
   fifo_reg_1_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n137, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_22_port);
   fifo_reg_1_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n139, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_21_port);
   fifo_reg_1_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n141, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_20_port);
   fifo_reg_1_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n143, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_19_port);
   fifo_reg_1_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n145, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_18_port);
   fifo_reg_1_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n147, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_17_port);
   fifo_reg_1_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n149, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_16_port);
   fifo_reg_1_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n151, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_15_port);
   fifo_reg_1_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n153, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_14_port);
   fifo_reg_1_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n155, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_13_port);
   fifo_reg_1_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n157, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_12_port);
   fifo_reg_1_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n159, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_11_port);
   fifo_reg_1_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n160, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_10_port);
   fifo_reg_1_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n161, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_9_port);
   fifo_reg_1_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n162, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_8_port);
   fifo_reg_1_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n163, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_7_port);
   fifo_reg_1_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n164, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_6_port);
   fifo_reg_1_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n165, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_5_port);
   fifo_reg_1_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n166, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_4_port);
   fifo_reg_0_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n231, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_3_port);
   fifo_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n232, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_2_port);
   fifo_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n233, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_1_port);
   fifo_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n234, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_0_port);
   fifo_reg_0_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n175, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_59_port);
   fifo_reg_0_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n176, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_58_port);
   fifo_reg_0_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n177, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_57_port);
   fifo_reg_0_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n178, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_56_port);
   fifo_reg_0_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n179, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_55_port);
   fifo_reg_0_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n180, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_54_port);
   fifo_reg_0_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n181, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_53_port);
   fifo_reg_0_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n182, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_52_port);
   fifo_reg_0_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n183, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_51_port);
   fifo_reg_0_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n184, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_50_port);
   fifo_reg_0_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n185, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_49_port);
   fifo_reg_0_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n186, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_48_port);
   fifo_reg_0_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n187, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_47_port);
   fifo_reg_0_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n188, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_46_port);
   fifo_reg_0_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n189, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_45_port);
   fifo_reg_0_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n190, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_44_port);
   fifo_reg_0_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n191, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_43_port);
   fifo_reg_0_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n192, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_42_port);
   fifo_reg_0_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n193, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_41_port);
   fifo_reg_0_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n194, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_40_port);
   fifo_reg_0_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n195, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_39_port);
   fifo_reg_0_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n196, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_38_port);
   fifo_reg_0_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n197, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_37_port);
   fifo_reg_0_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n198, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_36_port);
   fifo_reg_0_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n199, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_35_port);
   fifo_reg_0_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n200, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_34_port);
   fifo_reg_0_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n201, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_33_port);
   fifo_reg_0_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n202, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_32_port);
   fifo_reg_0_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n203, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_31_port);
   fifo_reg_0_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n204, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_30_port);
   fifo_reg_0_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n205, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_29_port);
   fifo_reg_0_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n206, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_28_port);
   fifo_reg_0_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n207, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_27_port);
   fifo_reg_0_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n208, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_26_port);
   fifo_reg_0_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n209, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_25_port);
   fifo_reg_0_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n210, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_24_port);
   fifo_reg_0_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n211, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_23_port);
   fifo_reg_0_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n212, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_22_port);
   fifo_reg_0_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n213, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_21_port);
   fifo_reg_0_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n214, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_20_port);
   fifo_reg_0_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n215, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_19_port);
   fifo_reg_0_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n216, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_18_port);
   fifo_reg_0_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n217, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_17_port);
   fifo_reg_0_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n218, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_16_port);
   fifo_reg_0_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n219, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_15_port);
   fifo_reg_0_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n220, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_14_port);
   fifo_reg_0_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n221, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_13_port);
   fifo_reg_0_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n222, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_12_port);
   fifo_reg_0_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n223, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_11_port);
   fifo_reg_0_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n224, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_10_port);
   fifo_reg_0_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n225, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_9_port);
   fifo_reg_0_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n226, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_8_port);
   fifo_reg_0_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n227, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_7_port);
   fifo_reg_0_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n228, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_6_port);
   fifo_reg_0_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n229, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_5_port);
   fifo_reg_0_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n230, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_4_port);
   valid_data_reg : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n235, CLK => clk, 
                           RESET => n47, SET => n1, QN => valid_data_port);
   read_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK 
                           => clk, RESET => n47, SET => n1, QN => 
                           read_pointer_0_port);
   U69 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U135 : INVx3_ASAP7_75t_R port map( A => rst, Y => n47);
   U138 : INVx1_ASAP7_75t_R port map( A => read_en, Y => n45);
   U140 : INVx1_ASAP7_75t_R port map( A => n29, Y => n17);
   U141 : INVx1_ASAP7_75t_R port map( A => n15, Y => n3);
   U142 : INVx1_ASAP7_75t_R port map( A => n31, Y => n43);
   U207 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n29);
   U208 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n15);
   U209 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n27);
   U210 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n25);
   U211 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n23);
   U212 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n21);
   U213 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n19);
   U214 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n13);
   U215 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n11);
   U216 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n9_port);
   U217 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n7_port);
   U218 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n5);
   U219 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n31);
   U220 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n33);
   U221 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n41);
   U222 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n39);
   U223 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n37);
   U224 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n35);
   U225 : INVx1_ASAP7_75t_R port map( A => N7, Y => N9);
   U226 : INVx1_ASAP7_75t_R port map( A => write_en, Y => n49);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity fifo_buff_depth2_10 is

   port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, clk, 
         rst : in std_logic;  data_out : out std_logic_vector (63 downto 0);  
         valid_data : out std_logic);

end fifo_buff_depth2_10;

architecture SYN_rtl of fifo_buff_depth2_10 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx3_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal valid_data_port, read_pointer_0_port, fifo_1_63_port, fifo_1_62_port,
      fifo_1_61_port, fifo_1_60_port, fifo_1_59_port, fifo_1_58_port, 
      fifo_1_57_port, fifo_1_56_port, fifo_1_55_port, fifo_1_54_port, 
      fifo_1_53_port, fifo_1_52_port, fifo_1_51_port, fifo_1_50_port, 
      fifo_1_49_port, fifo_1_48_port, fifo_1_47_port, fifo_1_46_port, 
      fifo_1_45_port, fifo_1_44_port, fifo_1_43_port, fifo_1_42_port, 
      fifo_1_41_port, fifo_1_40_port, fifo_1_39_port, fifo_1_38_port, 
      fifo_1_37_port, fifo_1_36_port, fifo_1_35_port, fifo_1_34_port, 
      fifo_1_33_port, fifo_1_32_port, fifo_1_31_port, fifo_1_30_port, 
      fifo_1_29_port, fifo_1_28_port, fifo_1_27_port, fifo_1_26_port, 
      fifo_1_25_port, fifo_1_24_port, fifo_1_23_port, fifo_1_22_port, 
      fifo_1_21_port, fifo_1_20_port, fifo_1_19_port, fifo_1_18_port, 
      fifo_1_17_port, fifo_1_16_port, fifo_1_15_port, fifo_1_14_port, 
      fifo_1_13_port, fifo_1_12_port, fifo_1_11_port, fifo_1_10_port, 
      fifo_1_9_port, fifo_1_8_port, fifo_1_7_port, fifo_1_6_port, fifo_1_5_port
      , fifo_1_4_port, fifo_1_3_port, fifo_1_2_port, fifo_1_1_port, 
      fifo_1_0_port, fifo_0_63_port, fifo_0_62_port, fifo_0_61_port, 
      fifo_0_60_port, fifo_0_59_port, fifo_0_58_port, fifo_0_57_port, 
      fifo_0_56_port, fifo_0_55_port, fifo_0_54_port, fifo_0_53_port, 
      fifo_0_52_port, fifo_0_51_port, fifo_0_50_port, fifo_0_49_port, 
      fifo_0_48_port, fifo_0_47_port, fifo_0_46_port, fifo_0_45_port, 
      fifo_0_44_port, fifo_0_43_port, fifo_0_42_port, fifo_0_41_port, 
      fifo_0_40_port, fifo_0_39_port, fifo_0_38_port, fifo_0_37_port, 
      fifo_0_36_port, fifo_0_35_port, fifo_0_34_port, fifo_0_33_port, 
      fifo_0_32_port, fifo_0_31_port, fifo_0_30_port, fifo_0_29_port, 
      fifo_0_28_port, fifo_0_27_port, fifo_0_26_port, fifo_0_25_port, 
      fifo_0_24_port, fifo_0_23_port, fifo_0_22_port, fifo_0_21_port, 
      fifo_0_20_port, fifo_0_19_port, fifo_0_18_port, fifo_0_17_port, 
      fifo_0_16_port, fifo_0_15_port, fifo_0_14_port, fifo_0_13_port, 
      fifo_0_12_port, fifo_0_11_port, fifo_0_10_port, fifo_0_9_port, 
      fifo_0_8_port, fifo_0_7_port, fifo_0_6_port, fifo_0_5_port, fifo_0_4_port
      , fifo_0_3_port, fifo_0_2_port, fifo_0_1_port, fifo_0_0_port, N7, N9, n1,
      n3, n5, n7_port, n9_port, n11, n13, n15, n17, n19, n21, n23, n25, n27, 
      n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57
      , n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, 
      n87, n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, n111, 
      n113, n115, n117, n119, n121, n123, n125, n127, n129, n131, n133, n135, 
      n137, n139, n141, n143, n145, n147, n149, n151, n153, n155, n157, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238 : std_logic;

begin
   valid_data <= valid_data_port;
   
   U4 : XOR2xp5_ASAP7_75t_R port map( A => N7, B => n43, Y => n238);
   U143 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_9_port, B1 => 
                           n43, B2 => fifo_0_9_port, Y => data_out(9));
   U144 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_8_port, B1 => 
                           n43, B2 => fifo_0_8_port, Y => data_out(8));
   U145 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_7_port, B1 => 
                           n43, B2 => fifo_0_7_port, Y => data_out(7));
   U146 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_6_port, B1 => 
                           n43, B2 => fifo_0_6_port, Y => data_out(6));
   U147 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_63_port, B1 => 
                           n43, B2 => fifo_0_63_port, Y => data_out(63));
   U148 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_62_port, B1 => 
                           n43, B2 => fifo_0_62_port, Y => data_out(62));
   U149 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_61_port, B1 => 
                           n43, B2 => fifo_0_61_port, Y => data_out(61));
   U150 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_60_port, B1 => 
                           n43, B2 => fifo_0_60_port, Y => data_out(60));
   U151 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_5_port, B1 => 
                           n43, B2 => fifo_0_5_port, Y => data_out(5));
   U152 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_59_port, B1 => 
                           n43, B2 => fifo_0_59_port, Y => data_out(59));
   U153 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_58_port, B1 => 
                           n43, B2 => fifo_0_58_port, Y => data_out(58));
   U154 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_57_port, B1 => 
                           n43, B2 => fifo_0_57_port, Y => data_out(57));
   U155 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_56_port, B1 => 
                           n43, B2 => fifo_0_56_port, Y => data_out(56));
   U156 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_55_port, B1 => 
                           n43, B2 => fifo_0_55_port, Y => data_out(55));
   U157 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_54_port, B1 => 
                           n43, B2 => fifo_0_54_port, Y => data_out(54));
   U158 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_53_port, B1 => 
                           n43, B2 => fifo_0_53_port, Y => data_out(53));
   U159 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_52_port, B1 => 
                           n43, B2 => fifo_0_52_port, Y => data_out(52));
   U160 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_51_port, B1 => 
                           n43, B2 => fifo_0_51_port, Y => data_out(51));
   U161 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_50_port, B1 => 
                           n43, B2 => fifo_0_50_port, Y => data_out(50));
   U162 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_4_port, B1 => 
                           n43, B2 => fifo_0_4_port, Y => data_out(4));
   U163 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_49_port, B1 => 
                           n43, B2 => fifo_0_49_port, Y => data_out(49));
   U164 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_48_port, B1 => 
                           n43, B2 => fifo_0_48_port, Y => data_out(48));
   U165 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_47_port, B1 => 
                           n43, B2 => fifo_0_47_port, Y => data_out(47));
   U166 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_46_port, B1 => 
                           n43, B2 => fifo_0_46_port, Y => data_out(46));
   U167 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_45_port, B1 => 
                           n43, B2 => fifo_0_45_port, Y => data_out(45));
   U168 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_44_port, B1 => 
                           n43, B2 => fifo_0_44_port, Y => data_out(44));
   U169 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_43_port, B1 => 
                           n43, B2 => fifo_0_43_port, Y => data_out(43));
   U170 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_42_port, B1 => 
                           n43, B2 => fifo_0_42_port, Y => data_out(42));
   U171 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_41_port, B1 => 
                           n43, B2 => fifo_0_41_port, Y => data_out(41));
   U172 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_40_port, B1 => 
                           n43, B2 => fifo_0_40_port, Y => data_out(40));
   U173 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_3_port, B1 => 
                           n43, B2 => fifo_0_3_port, Y => data_out(3));
   U174 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_39_port, B1 => 
                           n43, B2 => fifo_0_39_port, Y => data_out(39));
   U175 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_38_port, B1 => 
                           n43, B2 => fifo_0_38_port, Y => data_out(38));
   U176 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_37_port, B1 => 
                           n43, B2 => fifo_0_37_port, Y => data_out(37));
   U177 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_36_port, B1 => 
                           n43, B2 => fifo_0_36_port, Y => data_out(36));
   U178 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_35_port, B1 => 
                           n43, B2 => fifo_0_35_port, Y => data_out(35));
   U179 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_34_port, B1 => 
                           n43, B2 => fifo_0_34_port, Y => data_out(34));
   U180 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_33_port, B1 => 
                           n43, B2 => fifo_0_33_port, Y => data_out(33));
   U181 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_32_port, B1 => 
                           n43, B2 => fifo_0_32_port, Y => data_out(32));
   U182 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_31_port, B1 => 
                           n43, B2 => fifo_0_31_port, Y => data_out(31));
   U183 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_30_port, B1 => 
                           n43, B2 => fifo_0_30_port, Y => data_out(30));
   U184 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_2_port, B1 => 
                           n43, B2 => fifo_0_2_port, Y => data_out(2));
   U185 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_29_port, B1 => 
                           n43, B2 => fifo_0_29_port, Y => data_out(29));
   U186 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_28_port, B1 => 
                           n43, B2 => fifo_0_28_port, Y => data_out(28));
   U187 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_27_port, B1 => 
                           n43, B2 => fifo_0_27_port, Y => data_out(27));
   U188 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_26_port, B1 => 
                           n43, B2 => fifo_0_26_port, Y => data_out(26));
   U189 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_25_port, B1 => 
                           n43, B2 => fifo_0_25_port, Y => data_out(25));
   U190 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_24_port, B1 => 
                           n43, B2 => fifo_0_24_port, Y => data_out(24));
   U191 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_23_port, B1 => 
                           n43, B2 => fifo_0_23_port, Y => data_out(23));
   U192 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_22_port, B1 => 
                           n43, B2 => fifo_0_22_port, Y => data_out(22));
   U193 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_21_port, B1 => 
                           n43, B2 => fifo_0_21_port, Y => data_out(21));
   U194 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_20_port, B1 => 
                           n43, B2 => fifo_0_20_port, Y => data_out(20));
   U195 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_1_port, B1 => 
                           n43, B2 => fifo_0_1_port, Y => data_out(1));
   U196 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_19_port, B1 => 
                           n43, B2 => fifo_0_19_port, Y => data_out(19));
   U197 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_18_port, B1 => 
                           n43, B2 => fifo_0_18_port, Y => data_out(18));
   U198 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_17_port, B1 => 
                           n43, B2 => fifo_0_17_port, Y => data_out(17));
   U199 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_16_port, B1 => 
                           n43, B2 => fifo_0_16_port, Y => data_out(16));
   U200 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_15_port, B1 => 
                           n43, B2 => fifo_0_15_port, Y => data_out(15));
   U201 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_14_port, B1 => 
                           n43, B2 => fifo_0_14_port, Y => data_out(14));
   U202 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_13_port, B1 => 
                           n43, B2 => fifo_0_13_port, Y => data_out(13));
   U203 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_12_port, B1 => 
                           n43, B2 => fifo_0_12_port, Y => data_out(12));
   U204 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_11_port, B1 => 
                           n43, B2 => fifo_0_11_port, Y => data_out(11));
   U205 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_10_port, B1 => 
                           n43, B2 => fifo_0_10_port, Y => data_out(10));
   U206 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_0_port, B1 => 
                           n43, B2 => fifo_0_0_port, Y => data_out(0));
   U3 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n47, A2 => n238, B => 
                           valid_data_port, C => write_en, Y => n235);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_0_port, A2 => n17, B1 => 
                           data_in(0), B2 => n29, Y => n234);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_1_port, A2 => n17, B1 => 
                           data_in(1), B2 => n29, Y => n233);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_2_port, A2 => n17, B1 => 
                           data_in(2), B2 => n29, Y => n232);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_3_port, A2 => n17, B1 => 
                           data_in(3), B2 => n29, Y => n231);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_4_port, A2 => n17, B1 => 
                           data_in(4), B2 => n27, Y => n230);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_5_port, A2 => n17, B1 => 
                           data_in(5), B2 => n27, Y => n229);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_6_port, A2 => n17, B1 => 
                           data_in(6), B2 => n27, Y => n228);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_7_port, A2 => n17, B1 => 
                           data_in(7), B2 => n27, Y => n227);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_8_port, A2 => n17, B1 => 
                           data_in(8), B2 => n27, Y => n226);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_9_port, A2 => n17, B1 => 
                           data_in(9), B2 => n27, Y => n225);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_10_port, A2 => n17, B1 => 
                           data_in(10), B2 => n27, Y => n224);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_11_port, A2 => n17, B1 => 
                           data_in(11), B2 => n27, Y => n223);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_12_port, A2 => n17, B1 => 
                           data_in(12), B2 => n27, Y => n222);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_13_port, A2 => n17, B1 => 
                           data_in(13), B2 => n27, Y => n221);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_14_port, A2 => n17, B1 => 
                           data_in(14), B2 => n27, Y => n220);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_15_port, A2 => n17, B1 => 
                           data_in(15), B2 => n27, Y => n219);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_16_port, A2 => n17, B1 => 
                           data_in(16), B2 => n25, Y => n218);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_17_port, A2 => n17, B1 => 
                           data_in(17), B2 => n25, Y => n217);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_18_port, A2 => n17, B1 => 
                           data_in(18), B2 => n25, Y => n216);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_19_port, A2 => n17, B1 => 
                           data_in(19), B2 => n25, Y => n215);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_20_port, A2 => n17, B1 => 
                           data_in(20), B2 => n25, Y => n214);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_21_port, A2 => n17, B1 => 
                           data_in(21), B2 => n25, Y => n213);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_22_port, A2 => n17, B1 => 
                           data_in(22), B2 => n25, Y => n212);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_23_port, A2 => n17, B1 => 
                           data_in(23), B2 => n25, Y => n211);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_24_port, A2 => n17, B1 => 
                           data_in(24), B2 => n25, Y => n210);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_25_port, A2 => n17, B1 => 
                           data_in(25), B2 => n25, Y => n209);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_26_port, A2 => n17, B1 => 
                           data_in(26), B2 => n25, Y => n208);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_27_port, A2 => n17, B1 => 
                           data_in(27), B2 => n25, Y => n207);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_28_port, A2 => n17, B1 => 
                           data_in(28), B2 => n23, Y => n206);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_29_port, A2 => n17, B1 => 
                           data_in(29), B2 => n23, Y => n205);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_30_port, A2 => n17, B1 => 
                           data_in(30), B2 => n23, Y => n204);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_31_port, A2 => n17, B1 => 
                           data_in(31), B2 => n23, Y => n203);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_32_port, A2 => n17, B1 => 
                           data_in(32), B2 => n23, Y => n202);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_33_port, A2 => n17, B1 => 
                           data_in(33), B2 => n23, Y => n201);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_34_port, A2 => n17, B1 => 
                           data_in(34), B2 => n23, Y => n200);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_35_port, A2 => n17, B1 => 
                           data_in(35), B2 => n23, Y => n199);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_36_port, A2 => n17, B1 => 
                           data_in(36), B2 => n23, Y => n198);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_37_port, A2 => n17, B1 => 
                           data_in(37), B2 => n23, Y => n197);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_38_port, A2 => n17, B1 => 
                           data_in(38), B2 => n23, Y => n196);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_39_port, A2 => n17, B1 => 
                           data_in(39), B2 => n23, Y => n195);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_40_port, A2 => n17, B1 => 
                           data_in(40), B2 => n21, Y => n194);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_41_port, A2 => n17, B1 => 
                           data_in(41), B2 => n21, Y => n193);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_42_port, A2 => n17, B1 => 
                           data_in(42), B2 => n21, Y => n192);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_43_port, A2 => n17, B1 => 
                           data_in(43), B2 => n21, Y => n191);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_44_port, A2 => n17, B1 => 
                           data_in(44), B2 => n21, Y => n190);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_45_port, A2 => n17, B1 => 
                           data_in(45), B2 => n21, Y => n189);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_46_port, A2 => n17, B1 => 
                           data_in(46), B2 => n21, Y => n188);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_47_port, A2 => n17, B1 => 
                           data_in(47), B2 => n21, Y => n187);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_48_port, A2 => n17, B1 => 
                           data_in(48), B2 => n21, Y => n186);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_49_port, A2 => n17, B1 => 
                           data_in(49), B2 => n21, Y => n185);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_50_port, A2 => n17, B1 => 
                           data_in(50), B2 => n21, Y => n184);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_51_port, A2 => n17, B1 => 
                           data_in(51), B2 => n21, Y => n183);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_52_port, A2 => n17, B1 => 
                           data_in(52), B2 => n19, Y => n182);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_53_port, A2 => n17, B1 => 
                           data_in(53), B2 => n19, Y => n181);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_54_port, A2 => n17, B1 => 
                           data_in(54), B2 => n19, Y => n180);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_55_port, A2 => n17, B1 => 
                           data_in(55), B2 => n19, Y => n179);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_56_port, A2 => n17, B1 => 
                           data_in(56), B2 => n19, Y => n178);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_57_port, A2 => n17, B1 => 
                           data_in(57), B2 => n19, Y => n177);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_58_port, A2 => n17, B1 => 
                           data_in(58), B2 => n19, Y => n176);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_59_port, A2 => n17, B1 => 
                           data_in(59), B2 => n19, Y => n175);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_60_port, A2 => n17, B1 => 
                           data_in(60), B2 => n19, Y => n174);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_61_port, A2 => n17, B1 => 
                           data_in(61), B2 => n19, Y => n173);
   U67 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_62_port, A2 => n17, B1 => 
                           data_in(62), B2 => n19, Y => n172);
   U68 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_63_port, A2 => n17, B1 => 
                           data_in(63), B2 => n19, Y => n171);
   U70 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N9, Y => n237);
   U71 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_0_port, A2 => n3, B1 => 
                           data_in(0), B2 => n15, Y => n170);
   U72 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_1_port, A2 => n3, B1 => 
                           data_in(1), B2 => n15, Y => n169);
   U73 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_2_port, A2 => n3, B1 => 
                           data_in(2), B2 => n15, Y => n168);
   U74 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_3_port, A2 => n3, B1 => 
                           data_in(3), B2 => n15, Y => n167);
   U75 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_4_port, A2 => n3, B1 => 
                           data_in(4), B2 => n13, Y => n166);
   U76 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_5_port, A2 => n3, B1 => 
                           data_in(5), B2 => n13, Y => n165);
   U77 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_6_port, A2 => n3, B1 => 
                           data_in(6), B2 => n13, Y => n164);
   U78 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_7_port, A2 => n3, B1 => 
                           data_in(7), B2 => n13, Y => n163);
   U79 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_8_port, A2 => n3, B1 => 
                           data_in(8), B2 => n13, Y => n162);
   U80 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_9_port, A2 => n3, B1 => 
                           data_in(9), B2 => n13, Y => n161);
   U81 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_10_port, A2 => n3, B1 => 
                           data_in(10), B2 => n13, Y => n160);
   U82 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_11_port, A2 => n3, B1 => 
                           data_in(11), B2 => n13, Y => n159);
   U83 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_12_port, A2 => n3, B1 => 
                           data_in(12), B2 => n13, Y => n157);
   U84 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_13_port, A2 => n3, B1 => 
                           data_in(13), B2 => n13, Y => n155);
   U85 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_14_port, A2 => n3, B1 => 
                           data_in(14), B2 => n13, Y => n153);
   U86 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_15_port, A2 => n3, B1 => 
                           data_in(15), B2 => n13, Y => n151);
   U87 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_16_port, A2 => n3, B1 => 
                           data_in(16), B2 => n11, Y => n149);
   U88 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_17_port, A2 => n3, B1 => 
                           data_in(17), B2 => n11, Y => n147);
   U89 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_18_port, A2 => n3, B1 => 
                           data_in(18), B2 => n11, Y => n145);
   U90 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_19_port, A2 => n3, B1 => 
                           data_in(19), B2 => n11, Y => n143);
   U91 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_20_port, A2 => n3, B1 => 
                           data_in(20), B2 => n11, Y => n141);
   U92 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_21_port, A2 => n3, B1 => 
                           data_in(21), B2 => n11, Y => n139);
   U93 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_22_port, A2 => n3, B1 => 
                           data_in(22), B2 => n11, Y => n137);
   U94 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_23_port, A2 => n3, B1 => 
                           data_in(23), B2 => n11, Y => n135);
   U95 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_24_port, A2 => n3, B1 => 
                           data_in(24), B2 => n11, Y => n133);
   U96 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_25_port, A2 => n3, B1 => 
                           data_in(25), B2 => n11, Y => n131);
   U97 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_26_port, A2 => n3, B1 => 
                           data_in(26), B2 => n11, Y => n129);
   U98 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_27_port, A2 => n3, B1 => 
                           data_in(27), B2 => n11, Y => n127);
   U99 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_28_port, A2 => n3, B1 => 
                           data_in(28), B2 => n9_port, Y => n125);
   U100 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_29_port, A2 => n3, B1 => 
                           data_in(29), B2 => n9_port, Y => n123);
   U101 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_30_port, A2 => n3, B1 => 
                           data_in(30), B2 => n9_port, Y => n121);
   U102 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_31_port, A2 => n3, B1 => 
                           data_in(31), B2 => n9_port, Y => n119);
   U103 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_32_port, A2 => n3, B1 => 
                           data_in(32), B2 => n9_port, Y => n117);
   U104 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_33_port, A2 => n3, B1 => 
                           data_in(33), B2 => n9_port, Y => n115);
   U105 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_34_port, A2 => n3, B1 => 
                           data_in(34), B2 => n9_port, Y => n113);
   U106 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_35_port, A2 => n3, B1 => 
                           data_in(35), B2 => n9_port, Y => n111);
   U107 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_36_port, A2 => n3, B1 => 
                           data_in(36), B2 => n9_port, Y => n109);
   U108 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_37_port, A2 => n3, B1 => 
                           data_in(37), B2 => n9_port, Y => n107);
   U109 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_38_port, A2 => n3, B1 => 
                           data_in(38), B2 => n9_port, Y => n105);
   U110 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_39_port, A2 => n3, B1 => 
                           data_in(39), B2 => n9_port, Y => n103);
   U111 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_40_port, A2 => n3, B1 => 
                           data_in(40), B2 => n7_port, Y => n101);
   U112 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_41_port, A2 => n3, B1 => 
                           data_in(41), B2 => n7_port, Y => n99);
   U113 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_42_port, A2 => n3, B1 => 
                           data_in(42), B2 => n7_port, Y => n97);
   U114 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_43_port, A2 => n3, B1 => 
                           data_in(43), B2 => n7_port, Y => n95);
   U115 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_44_port, A2 => n3, B1 => 
                           data_in(44), B2 => n7_port, Y => n93);
   U116 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_45_port, A2 => n3, B1 => 
                           data_in(45), B2 => n7_port, Y => n91);
   U117 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_46_port, A2 => n3, B1 => 
                           data_in(46), B2 => n7_port, Y => n89);
   U118 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_47_port, A2 => n3, B1 => 
                           data_in(47), B2 => n7_port, Y => n87);
   U119 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_48_port, A2 => n3, B1 => 
                           data_in(48), B2 => n7_port, Y => n85);
   U120 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_49_port, A2 => n3, B1 => 
                           data_in(49), B2 => n7_port, Y => n83);
   U121 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_50_port, A2 => n3, B1 => 
                           data_in(50), B2 => n7_port, Y => n81);
   U122 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_51_port, A2 => n3, B1 => 
                           data_in(51), B2 => n7_port, Y => n79);
   U123 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_52_port, A2 => n3, B1 => 
                           data_in(52), B2 => n5, Y => n77);
   U124 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_53_port, A2 => n3, B1 => 
                           data_in(53), B2 => n5, Y => n75);
   U125 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_54_port, A2 => n3, B1 => 
                           data_in(54), B2 => n5, Y => n73);
   U126 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_55_port, A2 => n3, B1 => 
                           data_in(55), B2 => n5, Y => n71);
   U127 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_56_port, A2 => n3, B1 => 
                           data_in(56), B2 => n5, Y => n69);
   U128 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_57_port, A2 => n3, B1 => 
                           data_in(57), B2 => n5, Y => n67);
   U129 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_58_port, A2 => n3, B1 => 
                           data_in(58), B2 => n5, Y => n65);
   U130 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_59_port, A2 => n3, B1 => 
                           data_in(59), B2 => n5, Y => n63);
   U131 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_60_port, A2 => n3, B1 => 
                           data_in(60), B2 => n5, Y => n61);
   U132 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_61_port, A2 => n3, B1 => 
                           data_in(61), B2 => n5, Y => n59);
   U133 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_62_port, A2 => n3, B1 => 
                           data_in(62), B2 => n5, Y => n57);
   U134 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_63_port, A2 => n3, B1 => 
                           data_in(63), B2 => n5, Y => n55);
   U136 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N7, Y => n236);
   U137 : OAI22xp5_ASAP7_75t_R port map( A1 => n31, A2 => read_en, B1 => n43, 
                           B2 => n47, Y => n53);
   U139 : OAI22xp5_ASAP7_75t_R port map( A1 => N9, A2 => n49, B1 => write_en, 
                           B2 => N7, Y => n51);
   write_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK 
                           => clk, RESET => n45, SET => n1, QN => N7);
   fifo_reg_1_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n55, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_63_port);
   fifo_reg_1_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n57, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_62_port);
   fifo_reg_1_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n59, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_61_port);
   fifo_reg_1_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n61, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_60_port);
   fifo_reg_0_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n171, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_63_port);
   fifo_reg_0_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n172, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_62_port);
   fifo_reg_0_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n173, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_61_port);
   fifo_reg_0_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n174, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_60_port);
   fifo_reg_1_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n167, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_3_port);
   fifo_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n168, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_2_port);
   fifo_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n169, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_1_port);
   fifo_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n170, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_0_port);
   fifo_reg_1_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n63, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_59_port);
   fifo_reg_1_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n65, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_58_port);
   fifo_reg_1_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n67, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_57_port);
   fifo_reg_1_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n69, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_56_port);
   fifo_reg_1_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n71, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_55_port);
   fifo_reg_1_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n73, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_54_port);
   fifo_reg_1_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n75, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_53_port);
   fifo_reg_1_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n77, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_52_port);
   fifo_reg_1_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_51_port);
   fifo_reg_1_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_50_port);
   fifo_reg_1_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_49_port);
   fifo_reg_1_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_48_port);
   fifo_reg_1_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_47_port);
   fifo_reg_1_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_46_port);
   fifo_reg_1_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_45_port);
   fifo_reg_1_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_44_port);
   fifo_reg_1_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_43_port);
   fifo_reg_1_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_42_port);
   fifo_reg_1_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_41_port);
   fifo_reg_1_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_40_port);
   fifo_reg_1_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_39_port);
   fifo_reg_1_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_38_port);
   fifo_reg_1_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_37_port);
   fifo_reg_1_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_36_port);
   fifo_reg_1_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_35_port);
   fifo_reg_1_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_34_port);
   fifo_reg_1_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n115, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_33_port);
   fifo_reg_1_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n117, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_32_port);
   fifo_reg_1_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n119, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_31_port);
   fifo_reg_1_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n121, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_30_port);
   fifo_reg_1_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n123, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_29_port);
   fifo_reg_1_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n125, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_28_port);
   fifo_reg_1_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n127, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_27_port);
   fifo_reg_1_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n129, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_26_port);
   fifo_reg_1_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n131, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_25_port);
   fifo_reg_1_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n133, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_24_port);
   fifo_reg_1_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n135, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_23_port);
   fifo_reg_1_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n137, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_22_port);
   fifo_reg_1_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n139, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_21_port);
   fifo_reg_1_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n141, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_20_port);
   fifo_reg_1_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n143, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_19_port);
   fifo_reg_1_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n145, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_18_port);
   fifo_reg_1_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n147, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_17_port);
   fifo_reg_1_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n149, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_16_port);
   fifo_reg_1_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n151, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_15_port);
   fifo_reg_1_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n153, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_14_port);
   fifo_reg_1_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n155, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_13_port);
   fifo_reg_1_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n157, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_12_port);
   fifo_reg_1_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n159, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_11_port);
   fifo_reg_1_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n160, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_10_port);
   fifo_reg_1_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n161, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_9_port);
   fifo_reg_1_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n162, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_8_port);
   fifo_reg_1_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n163, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_7_port);
   fifo_reg_1_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n164, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_6_port);
   fifo_reg_1_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n165, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_5_port);
   fifo_reg_1_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n166, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_4_port);
   fifo_reg_0_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n231, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_3_port);
   fifo_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n232, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_2_port);
   fifo_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n233, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_1_port);
   fifo_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n234, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_0_port);
   fifo_reg_0_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n175, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_59_port);
   fifo_reg_0_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n176, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_58_port);
   fifo_reg_0_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n177, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_57_port);
   fifo_reg_0_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n178, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_56_port);
   fifo_reg_0_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n179, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_55_port);
   fifo_reg_0_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n180, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_54_port);
   fifo_reg_0_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n181, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_53_port);
   fifo_reg_0_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n182, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_52_port);
   fifo_reg_0_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n183, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_51_port);
   fifo_reg_0_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n184, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_50_port);
   fifo_reg_0_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n185, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_49_port);
   fifo_reg_0_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n186, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_48_port);
   fifo_reg_0_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n187, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_47_port);
   fifo_reg_0_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n188, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_46_port);
   fifo_reg_0_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n189, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_45_port);
   fifo_reg_0_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n190, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_44_port);
   fifo_reg_0_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n191, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_43_port);
   fifo_reg_0_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n192, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_42_port);
   fifo_reg_0_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n193, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_41_port);
   fifo_reg_0_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n194, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_40_port);
   fifo_reg_0_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n195, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_39_port);
   fifo_reg_0_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n196, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_38_port);
   fifo_reg_0_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n197, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_37_port);
   fifo_reg_0_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n198, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_36_port);
   fifo_reg_0_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n199, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_35_port);
   fifo_reg_0_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n200, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_34_port);
   fifo_reg_0_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n201, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_33_port);
   fifo_reg_0_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n202, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_32_port);
   fifo_reg_0_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n203, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_31_port);
   fifo_reg_0_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n204, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_30_port);
   fifo_reg_0_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n205, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_29_port);
   fifo_reg_0_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n206, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_28_port);
   fifo_reg_0_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n207, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_27_port);
   fifo_reg_0_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n208, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_26_port);
   fifo_reg_0_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n209, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_25_port);
   fifo_reg_0_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n210, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_24_port);
   fifo_reg_0_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n211, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_23_port);
   fifo_reg_0_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n212, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_22_port);
   fifo_reg_0_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n213, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_21_port);
   fifo_reg_0_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n214, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_20_port);
   fifo_reg_0_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n215, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_19_port);
   fifo_reg_0_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n216, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_18_port);
   fifo_reg_0_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n217, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_17_port);
   fifo_reg_0_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n218, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_16_port);
   fifo_reg_0_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n219, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_15_port);
   fifo_reg_0_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n220, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_14_port);
   fifo_reg_0_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n221, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_13_port);
   fifo_reg_0_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n222, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_12_port);
   fifo_reg_0_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n223, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_11_port);
   fifo_reg_0_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n224, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_10_port);
   fifo_reg_0_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n225, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_9_port);
   fifo_reg_0_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n226, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_8_port);
   fifo_reg_0_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n227, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_7_port);
   fifo_reg_0_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n228, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_6_port);
   fifo_reg_0_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n229, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_5_port);
   fifo_reg_0_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n230, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_4_port);
   valid_data_reg : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n235, CLK => clk, 
                           RESET => n45, SET => n1, QN => valid_data_port);
   read_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK 
                           => clk, RESET => n45, SET => n1, QN => 
                           read_pointer_0_port);
   U69 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U135 : INVx3_ASAP7_75t_R port map( A => rst, Y => n45);
   U138 : INVx1_ASAP7_75t_R port map( A => n29, Y => n17);
   U140 : INVx1_ASAP7_75t_R port map( A => n15, Y => n3);
   U141 : INVx1_ASAP7_75t_R port map( A => n31, Y => n43);
   U142 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n29);
   U207 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n15);
   U208 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n27);
   U209 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n25);
   U210 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n23);
   U211 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n21);
   U212 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n19);
   U213 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n13);
   U214 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n11);
   U215 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n9_port);
   U216 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n7_port);
   U217 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n5);
   U218 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n31);
   U219 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n33);
   U220 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n41);
   U221 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n39);
   U222 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n37);
   U223 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n35);
   U224 : INVx1_ASAP7_75t_R port map( A => read_en, Y => n47);
   U225 : INVx1_ASAP7_75t_R port map( A => N7, Y => N9);
   U226 : INVx1_ASAP7_75t_R port map( A => write_en, Y => n49);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity fifo_buff_depth2_9 is

   port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, clk, 
         rst : in std_logic;  data_out : out std_logic_vector (63 downto 0);  
         valid_data : out std_logic);

end fifo_buff_depth2_9;

architecture SYN_rtl of fifo_buff_depth2_9 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx3_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal valid_data_port, read_pointer_0_port, fifo_1_63_port, fifo_1_62_port,
      fifo_1_61_port, fifo_1_60_port, fifo_1_59_port, fifo_1_58_port, 
      fifo_1_57_port, fifo_1_56_port, fifo_1_55_port, fifo_1_54_port, 
      fifo_1_53_port, fifo_1_52_port, fifo_1_51_port, fifo_1_50_port, 
      fifo_1_49_port, fifo_1_48_port, fifo_1_47_port, fifo_1_46_port, 
      fifo_1_45_port, fifo_1_44_port, fifo_1_43_port, fifo_1_42_port, 
      fifo_1_41_port, fifo_1_40_port, fifo_1_39_port, fifo_1_38_port, 
      fifo_1_37_port, fifo_1_36_port, fifo_1_35_port, fifo_1_34_port, 
      fifo_1_33_port, fifo_1_32_port, fifo_1_31_port, fifo_1_30_port, 
      fifo_1_29_port, fifo_1_28_port, fifo_1_27_port, fifo_1_26_port, 
      fifo_1_25_port, fifo_1_24_port, fifo_1_23_port, fifo_1_22_port, 
      fifo_1_21_port, fifo_1_20_port, fifo_1_19_port, fifo_1_18_port, 
      fifo_1_17_port, fifo_1_16_port, fifo_1_15_port, fifo_1_14_port, 
      fifo_1_13_port, fifo_1_12_port, fifo_1_11_port, fifo_1_10_port, 
      fifo_1_9_port, fifo_1_8_port, fifo_1_7_port, fifo_1_6_port, fifo_1_5_port
      , fifo_1_4_port, fifo_1_3_port, fifo_1_2_port, fifo_1_1_port, 
      fifo_1_0_port, fifo_0_63_port, fifo_0_62_port, fifo_0_61_port, 
      fifo_0_60_port, fifo_0_59_port, fifo_0_58_port, fifo_0_57_port, 
      fifo_0_56_port, fifo_0_55_port, fifo_0_54_port, fifo_0_53_port, 
      fifo_0_52_port, fifo_0_51_port, fifo_0_50_port, fifo_0_49_port, 
      fifo_0_48_port, fifo_0_47_port, fifo_0_46_port, fifo_0_45_port, 
      fifo_0_44_port, fifo_0_43_port, fifo_0_42_port, fifo_0_41_port, 
      fifo_0_40_port, fifo_0_39_port, fifo_0_38_port, fifo_0_37_port, 
      fifo_0_36_port, fifo_0_35_port, fifo_0_34_port, fifo_0_33_port, 
      fifo_0_32_port, fifo_0_31_port, fifo_0_30_port, fifo_0_29_port, 
      fifo_0_28_port, fifo_0_27_port, fifo_0_26_port, fifo_0_25_port, 
      fifo_0_24_port, fifo_0_23_port, fifo_0_22_port, fifo_0_21_port, 
      fifo_0_20_port, fifo_0_19_port, fifo_0_18_port, fifo_0_17_port, 
      fifo_0_16_port, fifo_0_15_port, fifo_0_14_port, fifo_0_13_port, 
      fifo_0_12_port, fifo_0_11_port, fifo_0_10_port, fifo_0_9_port, 
      fifo_0_8_port, fifo_0_7_port, fifo_0_6_port, fifo_0_5_port, fifo_0_4_port
      , fifo_0_3_port, fifo_0_2_port, fifo_0_1_port, fifo_0_0_port, N7, N9, n1,
      n3, n5, n7_port, n9_port, n11, n13, n15, n17, n19, n21, n23, n25, n27, 
      n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57
      , n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, 
      n87, n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, n111, 
      n113, n115, n117, n119, n121, n123, n125, n127, n129, n131, n133, n135, 
      n137, n139, n141, n143, n145, n147, n149, n151, n153, n155, n157, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238 : std_logic;

begin
   valid_data <= valid_data_port;
   
   U4 : XOR2xp5_ASAP7_75t_R port map( A => N7, B => n43, Y => n238);
   U143 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_9_port, B1 => 
                           n43, B2 => fifo_0_9_port, Y => data_out(9));
   U144 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_8_port, B1 => 
                           n43, B2 => fifo_0_8_port, Y => data_out(8));
   U145 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_7_port, B1 => 
                           n43, B2 => fifo_0_7_port, Y => data_out(7));
   U146 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_6_port, B1 => 
                           n43, B2 => fifo_0_6_port, Y => data_out(6));
   U147 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_63_port, B1 => 
                           n43, B2 => fifo_0_63_port, Y => data_out(63));
   U148 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_62_port, B1 => 
                           n43, B2 => fifo_0_62_port, Y => data_out(62));
   U149 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_61_port, B1 => 
                           n43, B2 => fifo_0_61_port, Y => data_out(61));
   U150 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_60_port, B1 => 
                           n43, B2 => fifo_0_60_port, Y => data_out(60));
   U151 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_5_port, B1 => 
                           n43, B2 => fifo_0_5_port, Y => data_out(5));
   U152 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_59_port, B1 => 
                           n43, B2 => fifo_0_59_port, Y => data_out(59));
   U153 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_58_port, B1 => 
                           n43, B2 => fifo_0_58_port, Y => data_out(58));
   U154 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_57_port, B1 => 
                           n43, B2 => fifo_0_57_port, Y => data_out(57));
   U155 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_56_port, B1 => 
                           n43, B2 => fifo_0_56_port, Y => data_out(56));
   U156 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_55_port, B1 => 
                           n43, B2 => fifo_0_55_port, Y => data_out(55));
   U157 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_54_port, B1 => 
                           n43, B2 => fifo_0_54_port, Y => data_out(54));
   U158 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_53_port, B1 => 
                           n43, B2 => fifo_0_53_port, Y => data_out(53));
   U159 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_52_port, B1 => 
                           n43, B2 => fifo_0_52_port, Y => data_out(52));
   U160 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_51_port, B1 => 
                           n43, B2 => fifo_0_51_port, Y => data_out(51));
   U161 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_50_port, B1 => 
                           n43, B2 => fifo_0_50_port, Y => data_out(50));
   U162 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_4_port, B1 => 
                           n43, B2 => fifo_0_4_port, Y => data_out(4));
   U163 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_49_port, B1 => 
                           n43, B2 => fifo_0_49_port, Y => data_out(49));
   U164 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_48_port, B1 => 
                           n43, B2 => fifo_0_48_port, Y => data_out(48));
   U165 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_47_port, B1 => 
                           n43, B2 => fifo_0_47_port, Y => data_out(47));
   U166 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_46_port, B1 => 
                           n43, B2 => fifo_0_46_port, Y => data_out(46));
   U167 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_45_port, B1 => 
                           n43, B2 => fifo_0_45_port, Y => data_out(45));
   U168 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_44_port, B1 => 
                           n43, B2 => fifo_0_44_port, Y => data_out(44));
   U169 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_43_port, B1 => 
                           n43, B2 => fifo_0_43_port, Y => data_out(43));
   U170 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_42_port, B1 => 
                           n43, B2 => fifo_0_42_port, Y => data_out(42));
   U171 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_41_port, B1 => 
                           n43, B2 => fifo_0_41_port, Y => data_out(41));
   U172 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_40_port, B1 => 
                           n43, B2 => fifo_0_40_port, Y => data_out(40));
   U173 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_3_port, B1 => 
                           n43, B2 => fifo_0_3_port, Y => data_out(3));
   U174 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_39_port, B1 => 
                           n43, B2 => fifo_0_39_port, Y => data_out(39));
   U175 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_38_port, B1 => 
                           n43, B2 => fifo_0_38_port, Y => data_out(38));
   U176 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_37_port, B1 => 
                           n43, B2 => fifo_0_37_port, Y => data_out(37));
   U177 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_36_port, B1 => 
                           n43, B2 => fifo_0_36_port, Y => data_out(36));
   U178 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_35_port, B1 => 
                           n43, B2 => fifo_0_35_port, Y => data_out(35));
   U179 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_34_port, B1 => 
                           n43, B2 => fifo_0_34_port, Y => data_out(34));
   U180 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_33_port, B1 => 
                           n43, B2 => fifo_0_33_port, Y => data_out(33));
   U181 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_32_port, B1 => 
                           n43, B2 => fifo_0_32_port, Y => data_out(32));
   U182 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_31_port, B1 => 
                           n43, B2 => fifo_0_31_port, Y => data_out(31));
   U183 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_30_port, B1 => 
                           n43, B2 => fifo_0_30_port, Y => data_out(30));
   U184 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_2_port, B1 => 
                           n43, B2 => fifo_0_2_port, Y => data_out(2));
   U185 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_29_port, B1 => 
                           n43, B2 => fifo_0_29_port, Y => data_out(29));
   U186 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_28_port, B1 => 
                           n43, B2 => fifo_0_28_port, Y => data_out(28));
   U187 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_27_port, B1 => 
                           n43, B2 => fifo_0_27_port, Y => data_out(27));
   U188 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_26_port, B1 => 
                           n43, B2 => fifo_0_26_port, Y => data_out(26));
   U189 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_25_port, B1 => 
                           n43, B2 => fifo_0_25_port, Y => data_out(25));
   U190 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_24_port, B1 => 
                           n43, B2 => fifo_0_24_port, Y => data_out(24));
   U191 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_23_port, B1 => 
                           n43, B2 => fifo_0_23_port, Y => data_out(23));
   U192 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_22_port, B1 => 
                           n43, B2 => fifo_0_22_port, Y => data_out(22));
   U193 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_21_port, B1 => 
                           n43, B2 => fifo_0_21_port, Y => data_out(21));
   U194 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_20_port, B1 => 
                           n43, B2 => fifo_0_20_port, Y => data_out(20));
   U195 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_1_port, B1 => 
                           n43, B2 => fifo_0_1_port, Y => data_out(1));
   U196 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_19_port, B1 => 
                           n43, B2 => fifo_0_19_port, Y => data_out(19));
   U197 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_18_port, B1 => 
                           n43, B2 => fifo_0_18_port, Y => data_out(18));
   U198 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_17_port, B1 => 
                           n43, B2 => fifo_0_17_port, Y => data_out(17));
   U199 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_16_port, B1 => 
                           n43, B2 => fifo_0_16_port, Y => data_out(16));
   U200 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_15_port, B1 => 
                           n43, B2 => fifo_0_15_port, Y => data_out(15));
   U201 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_14_port, B1 => 
                           n43, B2 => fifo_0_14_port, Y => data_out(14));
   U202 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_13_port, B1 => 
                           n43, B2 => fifo_0_13_port, Y => data_out(13));
   U203 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_12_port, B1 => 
                           n43, B2 => fifo_0_12_port, Y => data_out(12));
   U204 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_11_port, B1 => 
                           n43, B2 => fifo_0_11_port, Y => data_out(11));
   U205 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_10_port, B1 => 
                           n43, B2 => fifo_0_10_port, Y => data_out(10));
   U206 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_0_port, B1 => 
                           n43, B2 => fifo_0_0_port, Y => data_out(0));
   U3 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n45, A2 => n238, B => 
                           valid_data_port, C => write_en, Y => n235);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_0_port, A2 => n17, B1 => 
                           data_in(0), B2 => n29, Y => n234);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_1_port, A2 => n17, B1 => 
                           data_in(1), B2 => n29, Y => n233);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_2_port, A2 => n17, B1 => 
                           data_in(2), B2 => n29, Y => n232);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_3_port, A2 => n17, B1 => 
                           data_in(3), B2 => n29, Y => n231);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_4_port, A2 => n17, B1 => 
                           data_in(4), B2 => n27, Y => n230);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_5_port, A2 => n17, B1 => 
                           data_in(5), B2 => n27, Y => n229);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_6_port, A2 => n17, B1 => 
                           data_in(6), B2 => n27, Y => n228);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_7_port, A2 => n17, B1 => 
                           data_in(7), B2 => n27, Y => n227);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_8_port, A2 => n17, B1 => 
                           data_in(8), B2 => n27, Y => n226);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_9_port, A2 => n17, B1 => 
                           data_in(9), B2 => n27, Y => n225);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_10_port, A2 => n17, B1 => 
                           data_in(10), B2 => n27, Y => n224);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_11_port, A2 => n17, B1 => 
                           data_in(11), B2 => n27, Y => n223);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_12_port, A2 => n17, B1 => 
                           data_in(12), B2 => n27, Y => n222);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_13_port, A2 => n17, B1 => 
                           data_in(13), B2 => n27, Y => n221);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_14_port, A2 => n17, B1 => 
                           data_in(14), B2 => n27, Y => n220);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_15_port, A2 => n17, B1 => 
                           data_in(15), B2 => n27, Y => n219);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_16_port, A2 => n17, B1 => 
                           data_in(16), B2 => n25, Y => n218);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_17_port, A2 => n17, B1 => 
                           data_in(17), B2 => n25, Y => n217);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_18_port, A2 => n17, B1 => 
                           data_in(18), B2 => n25, Y => n216);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_19_port, A2 => n17, B1 => 
                           data_in(19), B2 => n25, Y => n215);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_20_port, A2 => n17, B1 => 
                           data_in(20), B2 => n25, Y => n214);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_21_port, A2 => n17, B1 => 
                           data_in(21), B2 => n25, Y => n213);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_22_port, A2 => n17, B1 => 
                           data_in(22), B2 => n25, Y => n212);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_23_port, A2 => n17, B1 => 
                           data_in(23), B2 => n25, Y => n211);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_24_port, A2 => n17, B1 => 
                           data_in(24), B2 => n25, Y => n210);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_25_port, A2 => n17, B1 => 
                           data_in(25), B2 => n25, Y => n209);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_26_port, A2 => n17, B1 => 
                           data_in(26), B2 => n25, Y => n208);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_27_port, A2 => n17, B1 => 
                           data_in(27), B2 => n25, Y => n207);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_28_port, A2 => n17, B1 => 
                           data_in(28), B2 => n23, Y => n206);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_29_port, A2 => n17, B1 => 
                           data_in(29), B2 => n23, Y => n205);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_30_port, A2 => n17, B1 => 
                           data_in(30), B2 => n23, Y => n204);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_31_port, A2 => n17, B1 => 
                           data_in(31), B2 => n23, Y => n203);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_32_port, A2 => n17, B1 => 
                           data_in(32), B2 => n23, Y => n202);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_33_port, A2 => n17, B1 => 
                           data_in(33), B2 => n23, Y => n201);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_34_port, A2 => n17, B1 => 
                           data_in(34), B2 => n23, Y => n200);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_35_port, A2 => n17, B1 => 
                           data_in(35), B2 => n23, Y => n199);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_36_port, A2 => n17, B1 => 
                           data_in(36), B2 => n23, Y => n198);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_37_port, A2 => n17, B1 => 
                           data_in(37), B2 => n23, Y => n197);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_38_port, A2 => n17, B1 => 
                           data_in(38), B2 => n23, Y => n196);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_39_port, A2 => n17, B1 => 
                           data_in(39), B2 => n23, Y => n195);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_40_port, A2 => n17, B1 => 
                           data_in(40), B2 => n21, Y => n194);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_41_port, A2 => n17, B1 => 
                           data_in(41), B2 => n21, Y => n193);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_42_port, A2 => n17, B1 => 
                           data_in(42), B2 => n21, Y => n192);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_43_port, A2 => n17, B1 => 
                           data_in(43), B2 => n21, Y => n191);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_44_port, A2 => n17, B1 => 
                           data_in(44), B2 => n21, Y => n190);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_45_port, A2 => n17, B1 => 
                           data_in(45), B2 => n21, Y => n189);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_46_port, A2 => n17, B1 => 
                           data_in(46), B2 => n21, Y => n188);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_47_port, A2 => n17, B1 => 
                           data_in(47), B2 => n21, Y => n187);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_48_port, A2 => n17, B1 => 
                           data_in(48), B2 => n21, Y => n186);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_49_port, A2 => n17, B1 => 
                           data_in(49), B2 => n21, Y => n185);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_50_port, A2 => n17, B1 => 
                           data_in(50), B2 => n21, Y => n184);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_51_port, A2 => n17, B1 => 
                           data_in(51), B2 => n21, Y => n183);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_52_port, A2 => n17, B1 => 
                           data_in(52), B2 => n19, Y => n182);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_53_port, A2 => n17, B1 => 
                           data_in(53), B2 => n19, Y => n181);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_54_port, A2 => n17, B1 => 
                           data_in(54), B2 => n19, Y => n180);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_55_port, A2 => n17, B1 => 
                           data_in(55), B2 => n19, Y => n179);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_56_port, A2 => n17, B1 => 
                           data_in(56), B2 => n19, Y => n178);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_57_port, A2 => n17, B1 => 
                           data_in(57), B2 => n19, Y => n177);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_58_port, A2 => n17, B1 => 
                           data_in(58), B2 => n19, Y => n176);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_59_port, A2 => n17, B1 => 
                           data_in(59), B2 => n19, Y => n175);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_60_port, A2 => n17, B1 => 
                           data_in(60), B2 => n19, Y => n174);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_61_port, A2 => n17, B1 => 
                           data_in(61), B2 => n19, Y => n173);
   U67 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_62_port, A2 => n17, B1 => 
                           data_in(62), B2 => n19, Y => n172);
   U68 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_63_port, A2 => n17, B1 => 
                           data_in(63), B2 => n19, Y => n171);
   U70 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N9, Y => n237);
   U71 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_0_port, A2 => n3, B1 => 
                           data_in(0), B2 => n15, Y => n170);
   U72 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_1_port, A2 => n3, B1 => 
                           data_in(1), B2 => n15, Y => n169);
   U73 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_2_port, A2 => n3, B1 => 
                           data_in(2), B2 => n15, Y => n168);
   U74 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_3_port, A2 => n3, B1 => 
                           data_in(3), B2 => n15, Y => n167);
   U75 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_4_port, A2 => n3, B1 => 
                           data_in(4), B2 => n13, Y => n166);
   U76 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_5_port, A2 => n3, B1 => 
                           data_in(5), B2 => n13, Y => n165);
   U77 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_6_port, A2 => n3, B1 => 
                           data_in(6), B2 => n13, Y => n164);
   U78 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_7_port, A2 => n3, B1 => 
                           data_in(7), B2 => n13, Y => n163);
   U79 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_8_port, A2 => n3, B1 => 
                           data_in(8), B2 => n13, Y => n162);
   U80 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_9_port, A2 => n3, B1 => 
                           data_in(9), B2 => n13, Y => n161);
   U81 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_10_port, A2 => n3, B1 => 
                           data_in(10), B2 => n13, Y => n160);
   U82 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_11_port, A2 => n3, B1 => 
                           data_in(11), B2 => n13, Y => n159);
   U83 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_12_port, A2 => n3, B1 => 
                           data_in(12), B2 => n13, Y => n157);
   U84 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_13_port, A2 => n3, B1 => 
                           data_in(13), B2 => n13, Y => n155);
   U85 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_14_port, A2 => n3, B1 => 
                           data_in(14), B2 => n13, Y => n153);
   U86 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_15_port, A2 => n3, B1 => 
                           data_in(15), B2 => n13, Y => n151);
   U87 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_16_port, A2 => n3, B1 => 
                           data_in(16), B2 => n11, Y => n149);
   U88 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_17_port, A2 => n3, B1 => 
                           data_in(17), B2 => n11, Y => n147);
   U89 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_18_port, A2 => n3, B1 => 
                           data_in(18), B2 => n11, Y => n145);
   U90 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_19_port, A2 => n3, B1 => 
                           data_in(19), B2 => n11, Y => n143);
   U91 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_20_port, A2 => n3, B1 => 
                           data_in(20), B2 => n11, Y => n141);
   U92 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_21_port, A2 => n3, B1 => 
                           data_in(21), B2 => n11, Y => n139);
   U93 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_22_port, A2 => n3, B1 => 
                           data_in(22), B2 => n11, Y => n137);
   U94 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_23_port, A2 => n3, B1 => 
                           data_in(23), B2 => n11, Y => n135);
   U95 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_24_port, A2 => n3, B1 => 
                           data_in(24), B2 => n11, Y => n133);
   U96 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_25_port, A2 => n3, B1 => 
                           data_in(25), B2 => n11, Y => n131);
   U97 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_26_port, A2 => n3, B1 => 
                           data_in(26), B2 => n11, Y => n129);
   U98 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_27_port, A2 => n3, B1 => 
                           data_in(27), B2 => n11, Y => n127);
   U99 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_28_port, A2 => n3, B1 => 
                           data_in(28), B2 => n9_port, Y => n125);
   U100 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_29_port, A2 => n3, B1 => 
                           data_in(29), B2 => n9_port, Y => n123);
   U101 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_30_port, A2 => n3, B1 => 
                           data_in(30), B2 => n9_port, Y => n121);
   U102 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_31_port, A2 => n3, B1 => 
                           data_in(31), B2 => n9_port, Y => n119);
   U103 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_32_port, A2 => n3, B1 => 
                           data_in(32), B2 => n9_port, Y => n117);
   U104 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_33_port, A2 => n3, B1 => 
                           data_in(33), B2 => n9_port, Y => n115);
   U105 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_34_port, A2 => n3, B1 => 
                           data_in(34), B2 => n9_port, Y => n113);
   U106 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_35_port, A2 => n3, B1 => 
                           data_in(35), B2 => n9_port, Y => n111);
   U107 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_36_port, A2 => n3, B1 => 
                           data_in(36), B2 => n9_port, Y => n109);
   U108 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_37_port, A2 => n3, B1 => 
                           data_in(37), B2 => n9_port, Y => n107);
   U109 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_38_port, A2 => n3, B1 => 
                           data_in(38), B2 => n9_port, Y => n105);
   U110 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_39_port, A2 => n3, B1 => 
                           data_in(39), B2 => n9_port, Y => n103);
   U111 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_40_port, A2 => n3, B1 => 
                           data_in(40), B2 => n7_port, Y => n101);
   U112 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_41_port, A2 => n3, B1 => 
                           data_in(41), B2 => n7_port, Y => n99);
   U113 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_42_port, A2 => n3, B1 => 
                           data_in(42), B2 => n7_port, Y => n97);
   U114 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_43_port, A2 => n3, B1 => 
                           data_in(43), B2 => n7_port, Y => n95);
   U115 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_44_port, A2 => n3, B1 => 
                           data_in(44), B2 => n7_port, Y => n93);
   U116 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_45_port, A2 => n3, B1 => 
                           data_in(45), B2 => n7_port, Y => n91);
   U117 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_46_port, A2 => n3, B1 => 
                           data_in(46), B2 => n7_port, Y => n89);
   U118 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_47_port, A2 => n3, B1 => 
                           data_in(47), B2 => n7_port, Y => n87);
   U119 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_48_port, A2 => n3, B1 => 
                           data_in(48), B2 => n7_port, Y => n85);
   U120 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_49_port, A2 => n3, B1 => 
                           data_in(49), B2 => n7_port, Y => n83);
   U121 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_50_port, A2 => n3, B1 => 
                           data_in(50), B2 => n7_port, Y => n81);
   U122 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_51_port, A2 => n3, B1 => 
                           data_in(51), B2 => n7_port, Y => n79);
   U123 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_52_port, A2 => n3, B1 => 
                           data_in(52), B2 => n5, Y => n77);
   U124 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_53_port, A2 => n3, B1 => 
                           data_in(53), B2 => n5, Y => n75);
   U125 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_54_port, A2 => n3, B1 => 
                           data_in(54), B2 => n5, Y => n73);
   U126 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_55_port, A2 => n3, B1 => 
                           data_in(55), B2 => n5, Y => n71);
   U127 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_56_port, A2 => n3, B1 => 
                           data_in(56), B2 => n5, Y => n69);
   U128 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_57_port, A2 => n3, B1 => 
                           data_in(57), B2 => n5, Y => n67);
   U129 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_58_port, A2 => n3, B1 => 
                           data_in(58), B2 => n5, Y => n65);
   U130 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_59_port, A2 => n3, B1 => 
                           data_in(59), B2 => n5, Y => n63);
   U131 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_60_port, A2 => n3, B1 => 
                           data_in(60), B2 => n5, Y => n61);
   U132 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_61_port, A2 => n3, B1 => 
                           data_in(61), B2 => n5, Y => n59);
   U133 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_62_port, A2 => n3, B1 => 
                           data_in(62), B2 => n5, Y => n57);
   U134 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_63_port, A2 => n3, B1 => 
                           data_in(63), B2 => n5, Y => n55);
   U136 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N7, Y => n236);
   U137 : OAI22xp5_ASAP7_75t_R port map( A1 => n31, A2 => read_en, B1 => n43, 
                           B2 => n45, Y => n53);
   U139 : OAI22xp5_ASAP7_75t_R port map( A1 => N9, A2 => n49, B1 => write_en, 
                           B2 => N7, Y => n51);
   write_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK 
                           => clk, RESET => n47, SET => n1, QN => N7);
   fifo_reg_1_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n55, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_63_port);
   fifo_reg_1_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n57, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_62_port);
   fifo_reg_1_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n59, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_61_port);
   fifo_reg_1_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n61, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_60_port);
   fifo_reg_0_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n171, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_63_port);
   fifo_reg_0_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n172, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_62_port);
   fifo_reg_0_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n173, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_61_port);
   fifo_reg_0_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n174, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_60_port);
   fifo_reg_1_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n167, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_3_port);
   fifo_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n168, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_2_port);
   fifo_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n169, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_1_port);
   fifo_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n170, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_0_port);
   fifo_reg_1_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n63, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_59_port);
   fifo_reg_1_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n65, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_58_port);
   fifo_reg_1_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n67, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_57_port);
   fifo_reg_1_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n69, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_56_port);
   fifo_reg_1_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n71, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_55_port);
   fifo_reg_1_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n73, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_54_port);
   fifo_reg_1_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n75, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_53_port);
   fifo_reg_1_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n77, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_52_port);
   fifo_reg_1_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_51_port);
   fifo_reg_1_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_50_port);
   fifo_reg_1_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_49_port);
   fifo_reg_1_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_48_port);
   fifo_reg_1_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_47_port);
   fifo_reg_1_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_46_port);
   fifo_reg_1_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_45_port);
   fifo_reg_1_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_44_port);
   fifo_reg_1_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_43_port);
   fifo_reg_1_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_42_port);
   fifo_reg_1_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_41_port);
   fifo_reg_1_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_40_port);
   fifo_reg_1_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_39_port);
   fifo_reg_1_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_38_port);
   fifo_reg_1_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_37_port);
   fifo_reg_1_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_36_port);
   fifo_reg_1_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_35_port);
   fifo_reg_1_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_34_port);
   fifo_reg_1_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n115, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_33_port);
   fifo_reg_1_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n117, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_32_port);
   fifo_reg_1_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n119, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_31_port);
   fifo_reg_1_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n121, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_30_port);
   fifo_reg_1_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n123, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_29_port);
   fifo_reg_1_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n125, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_28_port);
   fifo_reg_1_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n127, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_27_port);
   fifo_reg_1_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n129, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_26_port);
   fifo_reg_1_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n131, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_25_port);
   fifo_reg_1_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n133, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_24_port);
   fifo_reg_1_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n135, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_23_port);
   fifo_reg_1_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n137, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_22_port);
   fifo_reg_1_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n139, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_21_port);
   fifo_reg_1_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n141, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_20_port);
   fifo_reg_1_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n143, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_19_port);
   fifo_reg_1_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n145, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_18_port);
   fifo_reg_1_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n147, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_17_port);
   fifo_reg_1_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n149, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_16_port);
   fifo_reg_1_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n151, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_15_port);
   fifo_reg_1_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n153, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_14_port);
   fifo_reg_1_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n155, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_13_port);
   fifo_reg_1_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n157, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_12_port);
   fifo_reg_1_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n159, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_11_port);
   fifo_reg_1_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n160, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_10_port);
   fifo_reg_1_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n161, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_9_port);
   fifo_reg_1_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n162, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_8_port);
   fifo_reg_1_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n163, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_7_port);
   fifo_reg_1_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n164, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_6_port);
   fifo_reg_1_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n165, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_5_port);
   fifo_reg_1_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n166, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_4_port);
   fifo_reg_0_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n231, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_3_port);
   fifo_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n232, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_2_port);
   fifo_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n233, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_1_port);
   fifo_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n234, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_0_port);
   fifo_reg_0_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n175, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_59_port);
   fifo_reg_0_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n176, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_58_port);
   fifo_reg_0_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n177, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_57_port);
   fifo_reg_0_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n178, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_56_port);
   fifo_reg_0_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n179, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_55_port);
   fifo_reg_0_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n180, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_54_port);
   fifo_reg_0_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n181, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_53_port);
   fifo_reg_0_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n182, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_52_port);
   fifo_reg_0_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n183, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_51_port);
   fifo_reg_0_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n184, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_50_port);
   fifo_reg_0_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n185, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_49_port);
   fifo_reg_0_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n186, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_48_port);
   fifo_reg_0_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n187, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_47_port);
   fifo_reg_0_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n188, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_46_port);
   fifo_reg_0_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n189, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_45_port);
   fifo_reg_0_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n190, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_44_port);
   fifo_reg_0_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n191, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_43_port);
   fifo_reg_0_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n192, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_42_port);
   fifo_reg_0_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n193, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_41_port);
   fifo_reg_0_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n194, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_40_port);
   fifo_reg_0_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n195, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_39_port);
   fifo_reg_0_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n196, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_38_port);
   fifo_reg_0_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n197, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_37_port);
   fifo_reg_0_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n198, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_36_port);
   fifo_reg_0_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n199, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_35_port);
   fifo_reg_0_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n200, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_34_port);
   fifo_reg_0_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n201, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_33_port);
   fifo_reg_0_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n202, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_32_port);
   fifo_reg_0_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n203, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_31_port);
   fifo_reg_0_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n204, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_30_port);
   fifo_reg_0_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n205, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_29_port);
   fifo_reg_0_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n206, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_28_port);
   fifo_reg_0_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n207, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_27_port);
   fifo_reg_0_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n208, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_26_port);
   fifo_reg_0_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n209, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_25_port);
   fifo_reg_0_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n210, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_24_port);
   fifo_reg_0_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n211, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_23_port);
   fifo_reg_0_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n212, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_22_port);
   fifo_reg_0_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n213, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_21_port);
   fifo_reg_0_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n214, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_20_port);
   fifo_reg_0_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n215, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_19_port);
   fifo_reg_0_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n216, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_18_port);
   fifo_reg_0_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n217, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_17_port);
   fifo_reg_0_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n218, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_16_port);
   fifo_reg_0_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n219, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_15_port);
   fifo_reg_0_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n220, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_14_port);
   fifo_reg_0_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n221, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_13_port);
   fifo_reg_0_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n222, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_12_port);
   fifo_reg_0_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n223, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_11_port);
   fifo_reg_0_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n224, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_10_port);
   fifo_reg_0_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n225, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_9_port);
   fifo_reg_0_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n226, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_8_port);
   fifo_reg_0_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n227, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_7_port);
   fifo_reg_0_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n228, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_6_port);
   fifo_reg_0_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n229, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_5_port);
   fifo_reg_0_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n230, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_4_port);
   valid_data_reg : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n235, CLK => clk, 
                           RESET => n47, SET => n1, QN => valid_data_port);
   read_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK 
                           => clk, RESET => n47, SET => n1, QN => 
                           read_pointer_0_port);
   U69 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U135 : INVx3_ASAP7_75t_R port map( A => rst, Y => n47);
   U138 : INVx1_ASAP7_75t_R port map( A => read_en, Y => n45);
   U140 : INVx1_ASAP7_75t_R port map( A => n29, Y => n17);
   U141 : INVx1_ASAP7_75t_R port map( A => n15, Y => n3);
   U142 : INVx1_ASAP7_75t_R port map( A => n31, Y => n43);
   U207 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n29);
   U208 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n15);
   U209 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n27);
   U210 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n25);
   U211 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n23);
   U212 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n21);
   U213 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n19);
   U214 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n13);
   U215 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n11);
   U216 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n9_port);
   U217 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n7_port);
   U218 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n5);
   U219 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n31);
   U220 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n33);
   U221 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n41);
   U222 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n39);
   U223 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n37);
   U224 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n35);
   U225 : INVx1_ASAP7_75t_R port map( A => N7, Y => N9);
   U226 : INVx1_ASAP7_75t_R port map( A => write_en, Y => n49);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity fifo_buff_depth2_8 is

   port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, clk, 
         rst : in std_logic;  data_out : out std_logic_vector (63 downto 0);  
         valid_data : out std_logic);

end fifo_buff_depth2_8;

architecture SYN_rtl of fifo_buff_depth2_8 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx3_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal valid_data_port, read_pointer_0_port, fifo_1_63_port, fifo_1_62_port,
      fifo_1_61_port, fifo_1_60_port, fifo_1_59_port, fifo_1_58_port, 
      fifo_1_57_port, fifo_1_56_port, fifo_1_55_port, fifo_1_54_port, 
      fifo_1_53_port, fifo_1_52_port, fifo_1_51_port, fifo_1_50_port, 
      fifo_1_49_port, fifo_1_48_port, fifo_1_47_port, fifo_1_46_port, 
      fifo_1_45_port, fifo_1_44_port, fifo_1_43_port, fifo_1_42_port, 
      fifo_1_41_port, fifo_1_40_port, fifo_1_39_port, fifo_1_38_port, 
      fifo_1_37_port, fifo_1_36_port, fifo_1_35_port, fifo_1_34_port, 
      fifo_1_33_port, fifo_1_32_port, fifo_1_31_port, fifo_1_30_port, 
      fifo_1_29_port, fifo_1_28_port, fifo_1_27_port, fifo_1_26_port, 
      fifo_1_25_port, fifo_1_24_port, fifo_1_23_port, fifo_1_22_port, 
      fifo_1_21_port, fifo_1_20_port, fifo_1_19_port, fifo_1_18_port, 
      fifo_1_17_port, fifo_1_16_port, fifo_1_15_port, fifo_1_14_port, 
      fifo_1_13_port, fifo_1_12_port, fifo_1_11_port, fifo_1_10_port, 
      fifo_1_9_port, fifo_1_8_port, fifo_1_7_port, fifo_1_6_port, fifo_1_5_port
      , fifo_1_4_port, fifo_1_3_port, fifo_1_2_port, fifo_1_1_port, 
      fifo_1_0_port, fifo_0_63_port, fifo_0_62_port, fifo_0_61_port, 
      fifo_0_60_port, fifo_0_59_port, fifo_0_58_port, fifo_0_57_port, 
      fifo_0_56_port, fifo_0_55_port, fifo_0_54_port, fifo_0_53_port, 
      fifo_0_52_port, fifo_0_51_port, fifo_0_50_port, fifo_0_49_port, 
      fifo_0_48_port, fifo_0_47_port, fifo_0_46_port, fifo_0_45_port, 
      fifo_0_44_port, fifo_0_43_port, fifo_0_42_port, fifo_0_41_port, 
      fifo_0_40_port, fifo_0_39_port, fifo_0_38_port, fifo_0_37_port, 
      fifo_0_36_port, fifo_0_35_port, fifo_0_34_port, fifo_0_33_port, 
      fifo_0_32_port, fifo_0_31_port, fifo_0_30_port, fifo_0_29_port, 
      fifo_0_28_port, fifo_0_27_port, fifo_0_26_port, fifo_0_25_port, 
      fifo_0_24_port, fifo_0_23_port, fifo_0_22_port, fifo_0_21_port, 
      fifo_0_20_port, fifo_0_19_port, fifo_0_18_port, fifo_0_17_port, 
      fifo_0_16_port, fifo_0_15_port, fifo_0_14_port, fifo_0_13_port, 
      fifo_0_12_port, fifo_0_11_port, fifo_0_10_port, fifo_0_9_port, 
      fifo_0_8_port, fifo_0_7_port, fifo_0_6_port, fifo_0_5_port, fifo_0_4_port
      , fifo_0_3_port, fifo_0_2_port, fifo_0_1_port, fifo_0_0_port, N7, N9, n1,
      n3, n5, n7_port, n9_port, n11, n13, n15, n17, n19, n21, n23, n25, n27, 
      n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57
      , n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, 
      n87, n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, n111, 
      n113, n115, n117, n119, n121, n123, n125, n127, n129, n131, n133, n135, 
      n137, n139, n141, n143, n145, n147, n149, n151, n153, n155, n157, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238 : std_logic;

begin
   valid_data <= valid_data_port;
   
   U4 : XOR2xp5_ASAP7_75t_R port map( A => N7, B => n43, Y => n238);
   U143 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_9_port, B1 => 
                           n43, B2 => fifo_0_9_port, Y => data_out(9));
   U144 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_8_port, B1 => 
                           n43, B2 => fifo_0_8_port, Y => data_out(8));
   U145 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_7_port, B1 => 
                           n43, B2 => fifo_0_7_port, Y => data_out(7));
   U146 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_6_port, B1 => 
                           n43, B2 => fifo_0_6_port, Y => data_out(6));
   U147 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_63_port, B1 => 
                           n43, B2 => fifo_0_63_port, Y => data_out(63));
   U148 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_62_port, B1 => 
                           n43, B2 => fifo_0_62_port, Y => data_out(62));
   U149 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_61_port, B1 => 
                           n43, B2 => fifo_0_61_port, Y => data_out(61));
   U150 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_60_port, B1 => 
                           n43, B2 => fifo_0_60_port, Y => data_out(60));
   U151 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_5_port, B1 => 
                           n43, B2 => fifo_0_5_port, Y => data_out(5));
   U152 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_59_port, B1 => 
                           n43, B2 => fifo_0_59_port, Y => data_out(59));
   U153 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_58_port, B1 => 
                           n43, B2 => fifo_0_58_port, Y => data_out(58));
   U154 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_57_port, B1 => 
                           n43, B2 => fifo_0_57_port, Y => data_out(57));
   U155 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_56_port, B1 => 
                           n43, B2 => fifo_0_56_port, Y => data_out(56));
   U156 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_55_port, B1 => 
                           n43, B2 => fifo_0_55_port, Y => data_out(55));
   U157 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_54_port, B1 => 
                           n43, B2 => fifo_0_54_port, Y => data_out(54));
   U158 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_53_port, B1 => 
                           n43, B2 => fifo_0_53_port, Y => data_out(53));
   U159 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_52_port, B1 => 
                           n43, B2 => fifo_0_52_port, Y => data_out(52));
   U160 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_51_port, B1 => 
                           n43, B2 => fifo_0_51_port, Y => data_out(51));
   U161 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_50_port, B1 => 
                           n43, B2 => fifo_0_50_port, Y => data_out(50));
   U162 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_4_port, B1 => 
                           n43, B2 => fifo_0_4_port, Y => data_out(4));
   U163 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_49_port, B1 => 
                           n43, B2 => fifo_0_49_port, Y => data_out(49));
   U164 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_48_port, B1 => 
                           n43, B2 => fifo_0_48_port, Y => data_out(48));
   U165 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_47_port, B1 => 
                           n43, B2 => fifo_0_47_port, Y => data_out(47));
   U166 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_46_port, B1 => 
                           n43, B2 => fifo_0_46_port, Y => data_out(46));
   U167 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_45_port, B1 => 
                           n43, B2 => fifo_0_45_port, Y => data_out(45));
   U168 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_44_port, B1 => 
                           n43, B2 => fifo_0_44_port, Y => data_out(44));
   U169 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_43_port, B1 => 
                           n43, B2 => fifo_0_43_port, Y => data_out(43));
   U170 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_42_port, B1 => 
                           n43, B2 => fifo_0_42_port, Y => data_out(42));
   U171 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_41_port, B1 => 
                           n43, B2 => fifo_0_41_port, Y => data_out(41));
   U172 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_40_port, B1 => 
                           n43, B2 => fifo_0_40_port, Y => data_out(40));
   U173 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_3_port, B1 => 
                           n43, B2 => fifo_0_3_port, Y => data_out(3));
   U174 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_39_port, B1 => 
                           n43, B2 => fifo_0_39_port, Y => data_out(39));
   U175 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_38_port, B1 => 
                           n43, B2 => fifo_0_38_port, Y => data_out(38));
   U176 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_37_port, B1 => 
                           n43, B2 => fifo_0_37_port, Y => data_out(37));
   U177 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_36_port, B1 => 
                           n43, B2 => fifo_0_36_port, Y => data_out(36));
   U178 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_35_port, B1 => 
                           n43, B2 => fifo_0_35_port, Y => data_out(35));
   U179 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_34_port, B1 => 
                           n43, B2 => fifo_0_34_port, Y => data_out(34));
   U180 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_33_port, B1 => 
                           n43, B2 => fifo_0_33_port, Y => data_out(33));
   U181 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_32_port, B1 => 
                           n43, B2 => fifo_0_32_port, Y => data_out(32));
   U182 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_31_port, B1 => 
                           n43, B2 => fifo_0_31_port, Y => data_out(31));
   U183 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_30_port, B1 => 
                           n43, B2 => fifo_0_30_port, Y => data_out(30));
   U184 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_2_port, B1 => 
                           n43, B2 => fifo_0_2_port, Y => data_out(2));
   U185 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_29_port, B1 => 
                           n43, B2 => fifo_0_29_port, Y => data_out(29));
   U186 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_28_port, B1 => 
                           n43, B2 => fifo_0_28_port, Y => data_out(28));
   U187 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_27_port, B1 => 
                           n43, B2 => fifo_0_27_port, Y => data_out(27));
   U188 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_26_port, B1 => 
                           n43, B2 => fifo_0_26_port, Y => data_out(26));
   U189 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_25_port, B1 => 
                           n43, B2 => fifo_0_25_port, Y => data_out(25));
   U190 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_24_port, B1 => 
                           n43, B2 => fifo_0_24_port, Y => data_out(24));
   U191 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_23_port, B1 => 
                           n43, B2 => fifo_0_23_port, Y => data_out(23));
   U192 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_22_port, B1 => 
                           n43, B2 => fifo_0_22_port, Y => data_out(22));
   U193 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_21_port, B1 => 
                           n43, B2 => fifo_0_21_port, Y => data_out(21));
   U194 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_20_port, B1 => 
                           n43, B2 => fifo_0_20_port, Y => data_out(20));
   U195 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_1_port, B1 => 
                           n43, B2 => fifo_0_1_port, Y => data_out(1));
   U196 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_19_port, B1 => 
                           n43, B2 => fifo_0_19_port, Y => data_out(19));
   U197 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_18_port, B1 => 
                           n43, B2 => fifo_0_18_port, Y => data_out(18));
   U198 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_17_port, B1 => 
                           n43, B2 => fifo_0_17_port, Y => data_out(17));
   U199 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_16_port, B1 => 
                           n43, B2 => fifo_0_16_port, Y => data_out(16));
   U200 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_15_port, B1 => 
                           n43, B2 => fifo_0_15_port, Y => data_out(15));
   U201 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_14_port, B1 => 
                           n43, B2 => fifo_0_14_port, Y => data_out(14));
   U202 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_13_port, B1 => 
                           n43, B2 => fifo_0_13_port, Y => data_out(13));
   U203 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_12_port, B1 => 
                           n43, B2 => fifo_0_12_port, Y => data_out(12));
   U204 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_11_port, B1 => 
                           n43, B2 => fifo_0_11_port, Y => data_out(11));
   U205 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_10_port, B1 => 
                           n43, B2 => fifo_0_10_port, Y => data_out(10));
   U206 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_0_port, B1 => 
                           n43, B2 => fifo_0_0_port, Y => data_out(0));
   U3 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n47, A2 => n238, B => 
                           valid_data_port, C => write_en, Y => n235);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_0_port, A2 => n17, B1 => 
                           data_in(0), B2 => n29, Y => n234);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_1_port, A2 => n17, B1 => 
                           data_in(1), B2 => n29, Y => n233);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_2_port, A2 => n17, B1 => 
                           data_in(2), B2 => n29, Y => n232);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_3_port, A2 => n17, B1 => 
                           data_in(3), B2 => n29, Y => n231);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_4_port, A2 => n17, B1 => 
                           data_in(4), B2 => n27, Y => n230);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_5_port, A2 => n17, B1 => 
                           data_in(5), B2 => n27, Y => n229);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_6_port, A2 => n17, B1 => 
                           data_in(6), B2 => n27, Y => n228);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_7_port, A2 => n17, B1 => 
                           data_in(7), B2 => n27, Y => n227);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_8_port, A2 => n17, B1 => 
                           data_in(8), B2 => n27, Y => n226);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_9_port, A2 => n17, B1 => 
                           data_in(9), B2 => n27, Y => n225);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_10_port, A2 => n17, B1 => 
                           data_in(10), B2 => n27, Y => n224);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_11_port, A2 => n17, B1 => 
                           data_in(11), B2 => n27, Y => n223);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_12_port, A2 => n17, B1 => 
                           data_in(12), B2 => n27, Y => n222);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_13_port, A2 => n17, B1 => 
                           data_in(13), B2 => n27, Y => n221);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_14_port, A2 => n17, B1 => 
                           data_in(14), B2 => n27, Y => n220);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_15_port, A2 => n17, B1 => 
                           data_in(15), B2 => n27, Y => n219);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_16_port, A2 => n17, B1 => 
                           data_in(16), B2 => n25, Y => n218);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_17_port, A2 => n17, B1 => 
                           data_in(17), B2 => n25, Y => n217);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_18_port, A2 => n17, B1 => 
                           data_in(18), B2 => n25, Y => n216);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_19_port, A2 => n17, B1 => 
                           data_in(19), B2 => n25, Y => n215);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_20_port, A2 => n17, B1 => 
                           data_in(20), B2 => n25, Y => n214);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_21_port, A2 => n17, B1 => 
                           data_in(21), B2 => n25, Y => n213);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_22_port, A2 => n17, B1 => 
                           data_in(22), B2 => n25, Y => n212);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_23_port, A2 => n17, B1 => 
                           data_in(23), B2 => n25, Y => n211);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_24_port, A2 => n17, B1 => 
                           data_in(24), B2 => n25, Y => n210);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_25_port, A2 => n17, B1 => 
                           data_in(25), B2 => n25, Y => n209);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_26_port, A2 => n17, B1 => 
                           data_in(26), B2 => n25, Y => n208);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_27_port, A2 => n17, B1 => 
                           data_in(27), B2 => n25, Y => n207);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_28_port, A2 => n17, B1 => 
                           data_in(28), B2 => n23, Y => n206);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_29_port, A2 => n17, B1 => 
                           data_in(29), B2 => n23, Y => n205);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_30_port, A2 => n17, B1 => 
                           data_in(30), B2 => n23, Y => n204);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_31_port, A2 => n17, B1 => 
                           data_in(31), B2 => n23, Y => n203);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_32_port, A2 => n17, B1 => 
                           data_in(32), B2 => n23, Y => n202);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_33_port, A2 => n17, B1 => 
                           data_in(33), B2 => n23, Y => n201);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_34_port, A2 => n17, B1 => 
                           data_in(34), B2 => n23, Y => n200);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_35_port, A2 => n17, B1 => 
                           data_in(35), B2 => n23, Y => n199);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_36_port, A2 => n17, B1 => 
                           data_in(36), B2 => n23, Y => n198);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_37_port, A2 => n17, B1 => 
                           data_in(37), B2 => n23, Y => n197);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_38_port, A2 => n17, B1 => 
                           data_in(38), B2 => n23, Y => n196);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_39_port, A2 => n17, B1 => 
                           data_in(39), B2 => n23, Y => n195);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_40_port, A2 => n17, B1 => 
                           data_in(40), B2 => n21, Y => n194);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_41_port, A2 => n17, B1 => 
                           data_in(41), B2 => n21, Y => n193);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_42_port, A2 => n17, B1 => 
                           data_in(42), B2 => n21, Y => n192);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_43_port, A2 => n17, B1 => 
                           data_in(43), B2 => n21, Y => n191);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_44_port, A2 => n17, B1 => 
                           data_in(44), B2 => n21, Y => n190);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_45_port, A2 => n17, B1 => 
                           data_in(45), B2 => n21, Y => n189);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_46_port, A2 => n17, B1 => 
                           data_in(46), B2 => n21, Y => n188);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_47_port, A2 => n17, B1 => 
                           data_in(47), B2 => n21, Y => n187);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_48_port, A2 => n17, B1 => 
                           data_in(48), B2 => n21, Y => n186);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_49_port, A2 => n17, B1 => 
                           data_in(49), B2 => n21, Y => n185);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_50_port, A2 => n17, B1 => 
                           data_in(50), B2 => n21, Y => n184);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_51_port, A2 => n17, B1 => 
                           data_in(51), B2 => n21, Y => n183);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_52_port, A2 => n17, B1 => 
                           data_in(52), B2 => n19, Y => n182);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_53_port, A2 => n17, B1 => 
                           data_in(53), B2 => n19, Y => n181);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_54_port, A2 => n17, B1 => 
                           data_in(54), B2 => n19, Y => n180);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_55_port, A2 => n17, B1 => 
                           data_in(55), B2 => n19, Y => n179);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_56_port, A2 => n17, B1 => 
                           data_in(56), B2 => n19, Y => n178);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_57_port, A2 => n17, B1 => 
                           data_in(57), B2 => n19, Y => n177);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_58_port, A2 => n17, B1 => 
                           data_in(58), B2 => n19, Y => n176);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_59_port, A2 => n17, B1 => 
                           data_in(59), B2 => n19, Y => n175);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_60_port, A2 => n17, B1 => 
                           data_in(60), B2 => n19, Y => n174);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_61_port, A2 => n17, B1 => 
                           data_in(61), B2 => n19, Y => n173);
   U67 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_62_port, A2 => n17, B1 => 
                           data_in(62), B2 => n19, Y => n172);
   U68 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_63_port, A2 => n17, B1 => 
                           data_in(63), B2 => n19, Y => n171);
   U70 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N9, Y => n237);
   U71 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_0_port, A2 => n3, B1 => 
                           data_in(0), B2 => n15, Y => n170);
   U72 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_1_port, A2 => n3, B1 => 
                           data_in(1), B2 => n15, Y => n169);
   U73 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_2_port, A2 => n3, B1 => 
                           data_in(2), B2 => n15, Y => n168);
   U74 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_3_port, A2 => n3, B1 => 
                           data_in(3), B2 => n15, Y => n167);
   U75 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_4_port, A2 => n3, B1 => 
                           data_in(4), B2 => n13, Y => n166);
   U76 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_5_port, A2 => n3, B1 => 
                           data_in(5), B2 => n13, Y => n165);
   U77 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_6_port, A2 => n3, B1 => 
                           data_in(6), B2 => n13, Y => n164);
   U78 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_7_port, A2 => n3, B1 => 
                           data_in(7), B2 => n13, Y => n163);
   U79 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_8_port, A2 => n3, B1 => 
                           data_in(8), B2 => n13, Y => n162);
   U80 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_9_port, A2 => n3, B1 => 
                           data_in(9), B2 => n13, Y => n161);
   U81 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_10_port, A2 => n3, B1 => 
                           data_in(10), B2 => n13, Y => n160);
   U82 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_11_port, A2 => n3, B1 => 
                           data_in(11), B2 => n13, Y => n159);
   U83 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_12_port, A2 => n3, B1 => 
                           data_in(12), B2 => n13, Y => n157);
   U84 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_13_port, A2 => n3, B1 => 
                           data_in(13), B2 => n13, Y => n155);
   U85 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_14_port, A2 => n3, B1 => 
                           data_in(14), B2 => n13, Y => n153);
   U86 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_15_port, A2 => n3, B1 => 
                           data_in(15), B2 => n13, Y => n151);
   U87 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_16_port, A2 => n3, B1 => 
                           data_in(16), B2 => n11, Y => n149);
   U88 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_17_port, A2 => n3, B1 => 
                           data_in(17), B2 => n11, Y => n147);
   U89 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_18_port, A2 => n3, B1 => 
                           data_in(18), B2 => n11, Y => n145);
   U90 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_19_port, A2 => n3, B1 => 
                           data_in(19), B2 => n11, Y => n143);
   U91 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_20_port, A2 => n3, B1 => 
                           data_in(20), B2 => n11, Y => n141);
   U92 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_21_port, A2 => n3, B1 => 
                           data_in(21), B2 => n11, Y => n139);
   U93 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_22_port, A2 => n3, B1 => 
                           data_in(22), B2 => n11, Y => n137);
   U94 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_23_port, A2 => n3, B1 => 
                           data_in(23), B2 => n11, Y => n135);
   U95 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_24_port, A2 => n3, B1 => 
                           data_in(24), B2 => n11, Y => n133);
   U96 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_25_port, A2 => n3, B1 => 
                           data_in(25), B2 => n11, Y => n131);
   U97 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_26_port, A2 => n3, B1 => 
                           data_in(26), B2 => n11, Y => n129);
   U98 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_27_port, A2 => n3, B1 => 
                           data_in(27), B2 => n11, Y => n127);
   U99 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_28_port, A2 => n3, B1 => 
                           data_in(28), B2 => n9_port, Y => n125);
   U100 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_29_port, A2 => n3, B1 => 
                           data_in(29), B2 => n9_port, Y => n123);
   U101 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_30_port, A2 => n3, B1 => 
                           data_in(30), B2 => n9_port, Y => n121);
   U102 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_31_port, A2 => n3, B1 => 
                           data_in(31), B2 => n9_port, Y => n119);
   U103 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_32_port, A2 => n3, B1 => 
                           data_in(32), B2 => n9_port, Y => n117);
   U104 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_33_port, A2 => n3, B1 => 
                           data_in(33), B2 => n9_port, Y => n115);
   U105 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_34_port, A2 => n3, B1 => 
                           data_in(34), B2 => n9_port, Y => n113);
   U106 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_35_port, A2 => n3, B1 => 
                           data_in(35), B2 => n9_port, Y => n111);
   U107 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_36_port, A2 => n3, B1 => 
                           data_in(36), B2 => n9_port, Y => n109);
   U108 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_37_port, A2 => n3, B1 => 
                           data_in(37), B2 => n9_port, Y => n107);
   U109 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_38_port, A2 => n3, B1 => 
                           data_in(38), B2 => n9_port, Y => n105);
   U110 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_39_port, A2 => n3, B1 => 
                           data_in(39), B2 => n9_port, Y => n103);
   U111 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_40_port, A2 => n3, B1 => 
                           data_in(40), B2 => n7_port, Y => n101);
   U112 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_41_port, A2 => n3, B1 => 
                           data_in(41), B2 => n7_port, Y => n99);
   U113 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_42_port, A2 => n3, B1 => 
                           data_in(42), B2 => n7_port, Y => n97);
   U114 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_43_port, A2 => n3, B1 => 
                           data_in(43), B2 => n7_port, Y => n95);
   U115 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_44_port, A2 => n3, B1 => 
                           data_in(44), B2 => n7_port, Y => n93);
   U116 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_45_port, A2 => n3, B1 => 
                           data_in(45), B2 => n7_port, Y => n91);
   U117 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_46_port, A2 => n3, B1 => 
                           data_in(46), B2 => n7_port, Y => n89);
   U118 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_47_port, A2 => n3, B1 => 
                           data_in(47), B2 => n7_port, Y => n87);
   U119 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_48_port, A2 => n3, B1 => 
                           data_in(48), B2 => n7_port, Y => n85);
   U120 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_49_port, A2 => n3, B1 => 
                           data_in(49), B2 => n7_port, Y => n83);
   U121 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_50_port, A2 => n3, B1 => 
                           data_in(50), B2 => n7_port, Y => n81);
   U122 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_51_port, A2 => n3, B1 => 
                           data_in(51), B2 => n7_port, Y => n79);
   U123 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_52_port, A2 => n3, B1 => 
                           data_in(52), B2 => n5, Y => n77);
   U124 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_53_port, A2 => n3, B1 => 
                           data_in(53), B2 => n5, Y => n75);
   U125 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_54_port, A2 => n3, B1 => 
                           data_in(54), B2 => n5, Y => n73);
   U126 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_55_port, A2 => n3, B1 => 
                           data_in(55), B2 => n5, Y => n71);
   U127 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_56_port, A2 => n3, B1 => 
                           data_in(56), B2 => n5, Y => n69);
   U128 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_57_port, A2 => n3, B1 => 
                           data_in(57), B2 => n5, Y => n67);
   U129 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_58_port, A2 => n3, B1 => 
                           data_in(58), B2 => n5, Y => n65);
   U130 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_59_port, A2 => n3, B1 => 
                           data_in(59), B2 => n5, Y => n63);
   U131 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_60_port, A2 => n3, B1 => 
                           data_in(60), B2 => n5, Y => n61);
   U132 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_61_port, A2 => n3, B1 => 
                           data_in(61), B2 => n5, Y => n59);
   U133 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_62_port, A2 => n3, B1 => 
                           data_in(62), B2 => n5, Y => n57);
   U134 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_63_port, A2 => n3, B1 => 
                           data_in(63), B2 => n5, Y => n55);
   U136 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N7, Y => n236);
   U137 : OAI22xp5_ASAP7_75t_R port map( A1 => n31, A2 => read_en, B1 => n43, 
                           B2 => n47, Y => n53);
   U139 : OAI22xp5_ASAP7_75t_R port map( A1 => N9, A2 => n49, B1 => write_en, 
                           B2 => N7, Y => n51);
   write_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK 
                           => clk, RESET => n45, SET => n1, QN => N7);
   fifo_reg_1_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n55, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_63_port);
   fifo_reg_1_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n57, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_62_port);
   fifo_reg_1_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n59, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_61_port);
   fifo_reg_1_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n61, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_60_port);
   fifo_reg_0_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n171, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_63_port);
   fifo_reg_0_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n172, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_62_port);
   fifo_reg_0_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n173, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_61_port);
   fifo_reg_0_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n174, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_60_port);
   fifo_reg_1_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n167, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_3_port);
   fifo_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n168, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_2_port);
   fifo_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n169, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_1_port);
   fifo_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n170, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_0_port);
   fifo_reg_1_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n63, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_59_port);
   fifo_reg_1_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n65, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_58_port);
   fifo_reg_1_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n67, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_57_port);
   fifo_reg_1_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n69, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_56_port);
   fifo_reg_1_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n71, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_55_port);
   fifo_reg_1_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n73, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_54_port);
   fifo_reg_1_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n75, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_53_port);
   fifo_reg_1_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n77, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_52_port);
   fifo_reg_1_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_51_port);
   fifo_reg_1_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_50_port);
   fifo_reg_1_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_49_port);
   fifo_reg_1_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_48_port);
   fifo_reg_1_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_47_port);
   fifo_reg_1_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_46_port);
   fifo_reg_1_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_45_port);
   fifo_reg_1_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_44_port);
   fifo_reg_1_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_43_port);
   fifo_reg_1_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_42_port);
   fifo_reg_1_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_41_port);
   fifo_reg_1_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_40_port);
   fifo_reg_1_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_39_port);
   fifo_reg_1_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_38_port);
   fifo_reg_1_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_37_port);
   fifo_reg_1_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_36_port);
   fifo_reg_1_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_35_port);
   fifo_reg_1_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_34_port);
   fifo_reg_1_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n115, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_33_port);
   fifo_reg_1_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n117, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_32_port);
   fifo_reg_1_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n119, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_31_port);
   fifo_reg_1_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n121, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_30_port);
   fifo_reg_1_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n123, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_29_port);
   fifo_reg_1_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n125, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_28_port);
   fifo_reg_1_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n127, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_27_port);
   fifo_reg_1_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n129, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_26_port);
   fifo_reg_1_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n131, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_25_port);
   fifo_reg_1_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n133, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_24_port);
   fifo_reg_1_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n135, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_23_port);
   fifo_reg_1_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n137, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_22_port);
   fifo_reg_1_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n139, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_21_port);
   fifo_reg_1_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n141, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_20_port);
   fifo_reg_1_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n143, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_19_port);
   fifo_reg_1_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n145, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_18_port);
   fifo_reg_1_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n147, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_17_port);
   fifo_reg_1_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n149, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_16_port);
   fifo_reg_1_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n151, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_15_port);
   fifo_reg_1_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n153, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_14_port);
   fifo_reg_1_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n155, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_13_port);
   fifo_reg_1_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n157, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_12_port);
   fifo_reg_1_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n159, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_11_port);
   fifo_reg_1_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n160, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_10_port);
   fifo_reg_1_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n161, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_9_port);
   fifo_reg_1_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n162, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_8_port);
   fifo_reg_1_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n163, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_7_port);
   fifo_reg_1_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n164, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_6_port);
   fifo_reg_1_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n165, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_5_port);
   fifo_reg_1_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n166, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_4_port);
   fifo_reg_0_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n231, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_3_port);
   fifo_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n232, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_2_port);
   fifo_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n233, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_1_port);
   fifo_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n234, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_0_port);
   fifo_reg_0_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n175, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_59_port);
   fifo_reg_0_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n176, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_58_port);
   fifo_reg_0_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n177, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_57_port);
   fifo_reg_0_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n178, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_56_port);
   fifo_reg_0_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n179, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_55_port);
   fifo_reg_0_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n180, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_54_port);
   fifo_reg_0_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n181, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_53_port);
   fifo_reg_0_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n182, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_52_port);
   fifo_reg_0_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n183, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_51_port);
   fifo_reg_0_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n184, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_50_port);
   fifo_reg_0_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n185, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_49_port);
   fifo_reg_0_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n186, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_48_port);
   fifo_reg_0_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n187, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_47_port);
   fifo_reg_0_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n188, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_46_port);
   fifo_reg_0_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n189, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_45_port);
   fifo_reg_0_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n190, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_44_port);
   fifo_reg_0_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n191, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_43_port);
   fifo_reg_0_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n192, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_42_port);
   fifo_reg_0_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n193, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_41_port);
   fifo_reg_0_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n194, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_40_port);
   fifo_reg_0_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n195, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_39_port);
   fifo_reg_0_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n196, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_38_port);
   fifo_reg_0_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n197, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_37_port);
   fifo_reg_0_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n198, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_36_port);
   fifo_reg_0_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n199, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_35_port);
   fifo_reg_0_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n200, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_34_port);
   fifo_reg_0_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n201, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_33_port);
   fifo_reg_0_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n202, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_32_port);
   fifo_reg_0_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n203, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_31_port);
   fifo_reg_0_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n204, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_30_port);
   fifo_reg_0_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n205, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_29_port);
   fifo_reg_0_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n206, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_28_port);
   fifo_reg_0_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n207, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_27_port);
   fifo_reg_0_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n208, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_26_port);
   fifo_reg_0_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n209, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_25_port);
   fifo_reg_0_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n210, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_24_port);
   fifo_reg_0_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n211, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_23_port);
   fifo_reg_0_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n212, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_22_port);
   fifo_reg_0_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n213, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_21_port);
   fifo_reg_0_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n214, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_20_port);
   fifo_reg_0_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n215, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_19_port);
   fifo_reg_0_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n216, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_18_port);
   fifo_reg_0_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n217, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_17_port);
   fifo_reg_0_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n218, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_16_port);
   fifo_reg_0_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n219, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_15_port);
   fifo_reg_0_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n220, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_14_port);
   fifo_reg_0_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n221, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_13_port);
   fifo_reg_0_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n222, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_12_port);
   fifo_reg_0_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n223, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_11_port);
   fifo_reg_0_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n224, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_10_port);
   fifo_reg_0_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n225, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_9_port);
   fifo_reg_0_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n226, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_8_port);
   fifo_reg_0_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n227, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_7_port);
   fifo_reg_0_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n228, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_6_port);
   fifo_reg_0_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n229, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_5_port);
   fifo_reg_0_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n230, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_4_port);
   valid_data_reg : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n235, CLK => clk, 
                           RESET => n45, SET => n1, QN => valid_data_port);
   read_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK 
                           => clk, RESET => n45, SET => n1, QN => 
                           read_pointer_0_port);
   U69 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U135 : INVx3_ASAP7_75t_R port map( A => rst, Y => n45);
   U138 : INVx1_ASAP7_75t_R port map( A => n29, Y => n17);
   U140 : INVx1_ASAP7_75t_R port map( A => n15, Y => n3);
   U141 : INVx1_ASAP7_75t_R port map( A => n31, Y => n43);
   U142 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n29);
   U207 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n15);
   U208 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n27);
   U209 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n25);
   U210 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n23);
   U211 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n21);
   U212 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n19);
   U213 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n13);
   U214 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n11);
   U215 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n9_port);
   U216 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n7_port);
   U217 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n5);
   U218 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n31);
   U219 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n33);
   U220 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n41);
   U221 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n39);
   U222 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n37);
   U223 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n35);
   U224 : INVx1_ASAP7_75t_R port map( A => read_en, Y => n47);
   U225 : INVx1_ASAP7_75t_R port map( A => N7, Y => N9);
   U226 : INVx1_ASAP7_75t_R port map( A => write_en, Y => n49);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity fifo_buff_depth2_7 is

   port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, clk, 
         rst : in std_logic;  data_out : out std_logic_vector (63 downto 0);  
         valid_data : out std_logic);

end fifo_buff_depth2_7;

architecture SYN_rtl of fifo_buff_depth2_7 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx3_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal valid_data_port, read_pointer_0_port, fifo_1_63_port, fifo_1_62_port,
      fifo_1_61_port, fifo_1_60_port, fifo_1_59_port, fifo_1_58_port, 
      fifo_1_57_port, fifo_1_56_port, fifo_1_55_port, fifo_1_54_port, 
      fifo_1_53_port, fifo_1_52_port, fifo_1_51_port, fifo_1_50_port, 
      fifo_1_49_port, fifo_1_48_port, fifo_1_47_port, fifo_1_46_port, 
      fifo_1_45_port, fifo_1_44_port, fifo_1_43_port, fifo_1_42_port, 
      fifo_1_41_port, fifo_1_40_port, fifo_1_39_port, fifo_1_38_port, 
      fifo_1_37_port, fifo_1_36_port, fifo_1_35_port, fifo_1_34_port, 
      fifo_1_33_port, fifo_1_32_port, fifo_1_31_port, fifo_1_30_port, 
      fifo_1_29_port, fifo_1_28_port, fifo_1_27_port, fifo_1_26_port, 
      fifo_1_25_port, fifo_1_24_port, fifo_1_23_port, fifo_1_22_port, 
      fifo_1_21_port, fifo_1_20_port, fifo_1_19_port, fifo_1_18_port, 
      fifo_1_17_port, fifo_1_16_port, fifo_1_15_port, fifo_1_14_port, 
      fifo_1_13_port, fifo_1_12_port, fifo_1_11_port, fifo_1_10_port, 
      fifo_1_9_port, fifo_1_8_port, fifo_1_7_port, fifo_1_6_port, fifo_1_5_port
      , fifo_1_4_port, fifo_1_3_port, fifo_1_2_port, fifo_1_1_port, 
      fifo_1_0_port, fifo_0_63_port, fifo_0_62_port, fifo_0_61_port, 
      fifo_0_60_port, fifo_0_59_port, fifo_0_58_port, fifo_0_57_port, 
      fifo_0_56_port, fifo_0_55_port, fifo_0_54_port, fifo_0_53_port, 
      fifo_0_52_port, fifo_0_51_port, fifo_0_50_port, fifo_0_49_port, 
      fifo_0_48_port, fifo_0_47_port, fifo_0_46_port, fifo_0_45_port, 
      fifo_0_44_port, fifo_0_43_port, fifo_0_42_port, fifo_0_41_port, 
      fifo_0_40_port, fifo_0_39_port, fifo_0_38_port, fifo_0_37_port, 
      fifo_0_36_port, fifo_0_35_port, fifo_0_34_port, fifo_0_33_port, 
      fifo_0_32_port, fifo_0_31_port, fifo_0_30_port, fifo_0_29_port, 
      fifo_0_28_port, fifo_0_27_port, fifo_0_26_port, fifo_0_25_port, 
      fifo_0_24_port, fifo_0_23_port, fifo_0_22_port, fifo_0_21_port, 
      fifo_0_20_port, fifo_0_19_port, fifo_0_18_port, fifo_0_17_port, 
      fifo_0_16_port, fifo_0_15_port, fifo_0_14_port, fifo_0_13_port, 
      fifo_0_12_port, fifo_0_11_port, fifo_0_10_port, fifo_0_9_port, 
      fifo_0_8_port, fifo_0_7_port, fifo_0_6_port, fifo_0_5_port, fifo_0_4_port
      , fifo_0_3_port, fifo_0_2_port, fifo_0_1_port, fifo_0_0_port, N7, N9, n1,
      n3, n5, n7_port, n9_port, n11, n13, n15, n17, n19, n21, n23, n25, n27, 
      n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57
      , n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, 
      n87, n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, n111, 
      n113, n115, n117, n119, n121, n123, n125, n127, n129, n131, n133, n135, 
      n137, n139, n141, n143, n145, n147, n149, n151, n153, n155, n157, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238 : std_logic;

begin
   valid_data <= valid_data_port;
   
   U4 : XOR2xp5_ASAP7_75t_R port map( A => N7, B => n43, Y => n238);
   U143 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_9_port, B1 => 
                           n43, B2 => fifo_0_9_port, Y => data_out(9));
   U144 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_8_port, B1 => 
                           n43, B2 => fifo_0_8_port, Y => data_out(8));
   U145 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_7_port, B1 => 
                           n43, B2 => fifo_0_7_port, Y => data_out(7));
   U146 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_6_port, B1 => 
                           n43, B2 => fifo_0_6_port, Y => data_out(6));
   U147 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_63_port, B1 => 
                           n43, B2 => fifo_0_63_port, Y => data_out(63));
   U148 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_62_port, B1 => 
                           n43, B2 => fifo_0_62_port, Y => data_out(62));
   U149 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_61_port, B1 => 
                           n43, B2 => fifo_0_61_port, Y => data_out(61));
   U150 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_60_port, B1 => 
                           n43, B2 => fifo_0_60_port, Y => data_out(60));
   U151 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_5_port, B1 => 
                           n43, B2 => fifo_0_5_port, Y => data_out(5));
   U152 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_59_port, B1 => 
                           n43, B2 => fifo_0_59_port, Y => data_out(59));
   U153 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_58_port, B1 => 
                           n43, B2 => fifo_0_58_port, Y => data_out(58));
   U154 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_57_port, B1 => 
                           n43, B2 => fifo_0_57_port, Y => data_out(57));
   U155 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_56_port, B1 => 
                           n43, B2 => fifo_0_56_port, Y => data_out(56));
   U156 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_55_port, B1 => 
                           n43, B2 => fifo_0_55_port, Y => data_out(55));
   U157 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_54_port, B1 => 
                           n43, B2 => fifo_0_54_port, Y => data_out(54));
   U158 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_53_port, B1 => 
                           n43, B2 => fifo_0_53_port, Y => data_out(53));
   U159 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_52_port, B1 => 
                           n43, B2 => fifo_0_52_port, Y => data_out(52));
   U160 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_51_port, B1 => 
                           n43, B2 => fifo_0_51_port, Y => data_out(51));
   U161 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_50_port, B1 => 
                           n43, B2 => fifo_0_50_port, Y => data_out(50));
   U162 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_4_port, B1 => 
                           n43, B2 => fifo_0_4_port, Y => data_out(4));
   U163 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_49_port, B1 => 
                           n43, B2 => fifo_0_49_port, Y => data_out(49));
   U164 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_48_port, B1 => 
                           n43, B2 => fifo_0_48_port, Y => data_out(48));
   U165 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_47_port, B1 => 
                           n43, B2 => fifo_0_47_port, Y => data_out(47));
   U166 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_46_port, B1 => 
                           n43, B2 => fifo_0_46_port, Y => data_out(46));
   U167 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_45_port, B1 => 
                           n43, B2 => fifo_0_45_port, Y => data_out(45));
   U168 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_44_port, B1 => 
                           n43, B2 => fifo_0_44_port, Y => data_out(44));
   U169 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_43_port, B1 => 
                           n43, B2 => fifo_0_43_port, Y => data_out(43));
   U170 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_42_port, B1 => 
                           n43, B2 => fifo_0_42_port, Y => data_out(42));
   U171 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_41_port, B1 => 
                           n43, B2 => fifo_0_41_port, Y => data_out(41));
   U172 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_40_port, B1 => 
                           n43, B2 => fifo_0_40_port, Y => data_out(40));
   U173 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_3_port, B1 => 
                           n43, B2 => fifo_0_3_port, Y => data_out(3));
   U174 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_39_port, B1 => 
                           n43, B2 => fifo_0_39_port, Y => data_out(39));
   U175 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_38_port, B1 => 
                           n43, B2 => fifo_0_38_port, Y => data_out(38));
   U176 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_37_port, B1 => 
                           n43, B2 => fifo_0_37_port, Y => data_out(37));
   U177 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_36_port, B1 => 
                           n43, B2 => fifo_0_36_port, Y => data_out(36));
   U178 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_35_port, B1 => 
                           n43, B2 => fifo_0_35_port, Y => data_out(35));
   U179 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_34_port, B1 => 
                           n43, B2 => fifo_0_34_port, Y => data_out(34));
   U180 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_33_port, B1 => 
                           n43, B2 => fifo_0_33_port, Y => data_out(33));
   U181 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_32_port, B1 => 
                           n43, B2 => fifo_0_32_port, Y => data_out(32));
   U182 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_31_port, B1 => 
                           n43, B2 => fifo_0_31_port, Y => data_out(31));
   U183 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_30_port, B1 => 
                           n43, B2 => fifo_0_30_port, Y => data_out(30));
   U184 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_2_port, B1 => 
                           n43, B2 => fifo_0_2_port, Y => data_out(2));
   U185 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_29_port, B1 => 
                           n43, B2 => fifo_0_29_port, Y => data_out(29));
   U186 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_28_port, B1 => 
                           n43, B2 => fifo_0_28_port, Y => data_out(28));
   U187 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_27_port, B1 => 
                           n43, B2 => fifo_0_27_port, Y => data_out(27));
   U188 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_26_port, B1 => 
                           n43, B2 => fifo_0_26_port, Y => data_out(26));
   U189 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_25_port, B1 => 
                           n43, B2 => fifo_0_25_port, Y => data_out(25));
   U190 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_24_port, B1 => 
                           n43, B2 => fifo_0_24_port, Y => data_out(24));
   U191 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_23_port, B1 => 
                           n43, B2 => fifo_0_23_port, Y => data_out(23));
   U192 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_22_port, B1 => 
                           n43, B2 => fifo_0_22_port, Y => data_out(22));
   U193 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_21_port, B1 => 
                           n43, B2 => fifo_0_21_port, Y => data_out(21));
   U194 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_20_port, B1 => 
                           n43, B2 => fifo_0_20_port, Y => data_out(20));
   U195 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_1_port, B1 => 
                           n43, B2 => fifo_0_1_port, Y => data_out(1));
   U196 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_19_port, B1 => 
                           n43, B2 => fifo_0_19_port, Y => data_out(19));
   U197 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_18_port, B1 => 
                           n43, B2 => fifo_0_18_port, Y => data_out(18));
   U198 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_17_port, B1 => 
                           n43, B2 => fifo_0_17_port, Y => data_out(17));
   U199 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_16_port, B1 => 
                           n43, B2 => fifo_0_16_port, Y => data_out(16));
   U200 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_15_port, B1 => 
                           n43, B2 => fifo_0_15_port, Y => data_out(15));
   U201 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_14_port, B1 => 
                           n43, B2 => fifo_0_14_port, Y => data_out(14));
   U202 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_13_port, B1 => 
                           n43, B2 => fifo_0_13_port, Y => data_out(13));
   U203 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_12_port, B1 => 
                           n43, B2 => fifo_0_12_port, Y => data_out(12));
   U204 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_11_port, B1 => 
                           n43, B2 => fifo_0_11_port, Y => data_out(11));
   U205 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_10_port, B1 => 
                           n43, B2 => fifo_0_10_port, Y => data_out(10));
   U206 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_0_port, B1 => 
                           n43, B2 => fifo_0_0_port, Y => data_out(0));
   U3 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n45, A2 => n238, B => 
                           valid_data_port, C => write_en, Y => n235);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_0_port, A2 => n17, B1 => 
                           data_in(0), B2 => n29, Y => n234);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_1_port, A2 => n17, B1 => 
                           data_in(1), B2 => n29, Y => n233);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_2_port, A2 => n17, B1 => 
                           data_in(2), B2 => n29, Y => n232);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_3_port, A2 => n17, B1 => 
                           data_in(3), B2 => n29, Y => n231);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_4_port, A2 => n17, B1 => 
                           data_in(4), B2 => n27, Y => n230);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_5_port, A2 => n17, B1 => 
                           data_in(5), B2 => n27, Y => n229);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_6_port, A2 => n17, B1 => 
                           data_in(6), B2 => n27, Y => n228);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_7_port, A2 => n17, B1 => 
                           data_in(7), B2 => n27, Y => n227);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_8_port, A2 => n17, B1 => 
                           data_in(8), B2 => n27, Y => n226);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_9_port, A2 => n17, B1 => 
                           data_in(9), B2 => n27, Y => n225);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_10_port, A2 => n17, B1 => 
                           data_in(10), B2 => n27, Y => n224);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_11_port, A2 => n17, B1 => 
                           data_in(11), B2 => n27, Y => n223);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_12_port, A2 => n17, B1 => 
                           data_in(12), B2 => n27, Y => n222);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_13_port, A2 => n17, B1 => 
                           data_in(13), B2 => n27, Y => n221);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_14_port, A2 => n17, B1 => 
                           data_in(14), B2 => n27, Y => n220);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_15_port, A2 => n17, B1 => 
                           data_in(15), B2 => n27, Y => n219);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_16_port, A2 => n17, B1 => 
                           data_in(16), B2 => n25, Y => n218);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_17_port, A2 => n17, B1 => 
                           data_in(17), B2 => n25, Y => n217);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_18_port, A2 => n17, B1 => 
                           data_in(18), B2 => n25, Y => n216);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_19_port, A2 => n17, B1 => 
                           data_in(19), B2 => n25, Y => n215);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_20_port, A2 => n17, B1 => 
                           data_in(20), B2 => n25, Y => n214);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_21_port, A2 => n17, B1 => 
                           data_in(21), B2 => n25, Y => n213);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_22_port, A2 => n17, B1 => 
                           data_in(22), B2 => n25, Y => n212);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_23_port, A2 => n17, B1 => 
                           data_in(23), B2 => n25, Y => n211);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_24_port, A2 => n17, B1 => 
                           data_in(24), B2 => n25, Y => n210);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_25_port, A2 => n17, B1 => 
                           data_in(25), B2 => n25, Y => n209);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_26_port, A2 => n17, B1 => 
                           data_in(26), B2 => n25, Y => n208);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_27_port, A2 => n17, B1 => 
                           data_in(27), B2 => n25, Y => n207);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_28_port, A2 => n17, B1 => 
                           data_in(28), B2 => n23, Y => n206);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_29_port, A2 => n17, B1 => 
                           data_in(29), B2 => n23, Y => n205);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_30_port, A2 => n17, B1 => 
                           data_in(30), B2 => n23, Y => n204);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_31_port, A2 => n17, B1 => 
                           data_in(31), B2 => n23, Y => n203);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_32_port, A2 => n17, B1 => 
                           data_in(32), B2 => n23, Y => n202);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_33_port, A2 => n17, B1 => 
                           data_in(33), B2 => n23, Y => n201);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_34_port, A2 => n17, B1 => 
                           data_in(34), B2 => n23, Y => n200);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_35_port, A2 => n17, B1 => 
                           data_in(35), B2 => n23, Y => n199);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_36_port, A2 => n17, B1 => 
                           data_in(36), B2 => n23, Y => n198);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_37_port, A2 => n17, B1 => 
                           data_in(37), B2 => n23, Y => n197);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_38_port, A2 => n17, B1 => 
                           data_in(38), B2 => n23, Y => n196);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_39_port, A2 => n17, B1 => 
                           data_in(39), B2 => n23, Y => n195);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_40_port, A2 => n17, B1 => 
                           data_in(40), B2 => n21, Y => n194);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_41_port, A2 => n17, B1 => 
                           data_in(41), B2 => n21, Y => n193);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_42_port, A2 => n17, B1 => 
                           data_in(42), B2 => n21, Y => n192);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_43_port, A2 => n17, B1 => 
                           data_in(43), B2 => n21, Y => n191);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_44_port, A2 => n17, B1 => 
                           data_in(44), B2 => n21, Y => n190);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_45_port, A2 => n17, B1 => 
                           data_in(45), B2 => n21, Y => n189);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_46_port, A2 => n17, B1 => 
                           data_in(46), B2 => n21, Y => n188);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_47_port, A2 => n17, B1 => 
                           data_in(47), B2 => n21, Y => n187);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_48_port, A2 => n17, B1 => 
                           data_in(48), B2 => n21, Y => n186);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_49_port, A2 => n17, B1 => 
                           data_in(49), B2 => n21, Y => n185);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_50_port, A2 => n17, B1 => 
                           data_in(50), B2 => n21, Y => n184);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_51_port, A2 => n17, B1 => 
                           data_in(51), B2 => n21, Y => n183);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_52_port, A2 => n17, B1 => 
                           data_in(52), B2 => n19, Y => n182);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_53_port, A2 => n17, B1 => 
                           data_in(53), B2 => n19, Y => n181);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_54_port, A2 => n17, B1 => 
                           data_in(54), B2 => n19, Y => n180);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_55_port, A2 => n17, B1 => 
                           data_in(55), B2 => n19, Y => n179);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_56_port, A2 => n17, B1 => 
                           data_in(56), B2 => n19, Y => n178);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_57_port, A2 => n17, B1 => 
                           data_in(57), B2 => n19, Y => n177);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_58_port, A2 => n17, B1 => 
                           data_in(58), B2 => n19, Y => n176);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_59_port, A2 => n17, B1 => 
                           data_in(59), B2 => n19, Y => n175);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_60_port, A2 => n17, B1 => 
                           data_in(60), B2 => n19, Y => n174);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_61_port, A2 => n17, B1 => 
                           data_in(61), B2 => n19, Y => n173);
   U67 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_62_port, A2 => n17, B1 => 
                           data_in(62), B2 => n19, Y => n172);
   U68 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_63_port, A2 => n17, B1 => 
                           data_in(63), B2 => n19, Y => n171);
   U70 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N9, Y => n237);
   U71 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_0_port, A2 => n3, B1 => 
                           data_in(0), B2 => n15, Y => n170);
   U72 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_1_port, A2 => n3, B1 => 
                           data_in(1), B2 => n15, Y => n169);
   U73 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_2_port, A2 => n3, B1 => 
                           data_in(2), B2 => n15, Y => n168);
   U74 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_3_port, A2 => n3, B1 => 
                           data_in(3), B2 => n15, Y => n167);
   U75 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_4_port, A2 => n3, B1 => 
                           data_in(4), B2 => n13, Y => n166);
   U76 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_5_port, A2 => n3, B1 => 
                           data_in(5), B2 => n13, Y => n165);
   U77 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_6_port, A2 => n3, B1 => 
                           data_in(6), B2 => n13, Y => n164);
   U78 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_7_port, A2 => n3, B1 => 
                           data_in(7), B2 => n13, Y => n163);
   U79 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_8_port, A2 => n3, B1 => 
                           data_in(8), B2 => n13, Y => n162);
   U80 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_9_port, A2 => n3, B1 => 
                           data_in(9), B2 => n13, Y => n161);
   U81 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_10_port, A2 => n3, B1 => 
                           data_in(10), B2 => n13, Y => n160);
   U82 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_11_port, A2 => n3, B1 => 
                           data_in(11), B2 => n13, Y => n159);
   U83 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_12_port, A2 => n3, B1 => 
                           data_in(12), B2 => n13, Y => n157);
   U84 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_13_port, A2 => n3, B1 => 
                           data_in(13), B2 => n13, Y => n155);
   U85 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_14_port, A2 => n3, B1 => 
                           data_in(14), B2 => n13, Y => n153);
   U86 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_15_port, A2 => n3, B1 => 
                           data_in(15), B2 => n13, Y => n151);
   U87 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_16_port, A2 => n3, B1 => 
                           data_in(16), B2 => n11, Y => n149);
   U88 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_17_port, A2 => n3, B1 => 
                           data_in(17), B2 => n11, Y => n147);
   U89 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_18_port, A2 => n3, B1 => 
                           data_in(18), B2 => n11, Y => n145);
   U90 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_19_port, A2 => n3, B1 => 
                           data_in(19), B2 => n11, Y => n143);
   U91 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_20_port, A2 => n3, B1 => 
                           data_in(20), B2 => n11, Y => n141);
   U92 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_21_port, A2 => n3, B1 => 
                           data_in(21), B2 => n11, Y => n139);
   U93 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_22_port, A2 => n3, B1 => 
                           data_in(22), B2 => n11, Y => n137);
   U94 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_23_port, A2 => n3, B1 => 
                           data_in(23), B2 => n11, Y => n135);
   U95 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_24_port, A2 => n3, B1 => 
                           data_in(24), B2 => n11, Y => n133);
   U96 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_25_port, A2 => n3, B1 => 
                           data_in(25), B2 => n11, Y => n131);
   U97 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_26_port, A2 => n3, B1 => 
                           data_in(26), B2 => n11, Y => n129);
   U98 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_27_port, A2 => n3, B1 => 
                           data_in(27), B2 => n11, Y => n127);
   U99 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_28_port, A2 => n3, B1 => 
                           data_in(28), B2 => n9_port, Y => n125);
   U100 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_29_port, A2 => n3, B1 => 
                           data_in(29), B2 => n9_port, Y => n123);
   U101 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_30_port, A2 => n3, B1 => 
                           data_in(30), B2 => n9_port, Y => n121);
   U102 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_31_port, A2 => n3, B1 => 
                           data_in(31), B2 => n9_port, Y => n119);
   U103 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_32_port, A2 => n3, B1 => 
                           data_in(32), B2 => n9_port, Y => n117);
   U104 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_33_port, A2 => n3, B1 => 
                           data_in(33), B2 => n9_port, Y => n115);
   U105 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_34_port, A2 => n3, B1 => 
                           data_in(34), B2 => n9_port, Y => n113);
   U106 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_35_port, A2 => n3, B1 => 
                           data_in(35), B2 => n9_port, Y => n111);
   U107 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_36_port, A2 => n3, B1 => 
                           data_in(36), B2 => n9_port, Y => n109);
   U108 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_37_port, A2 => n3, B1 => 
                           data_in(37), B2 => n9_port, Y => n107);
   U109 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_38_port, A2 => n3, B1 => 
                           data_in(38), B2 => n9_port, Y => n105);
   U110 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_39_port, A2 => n3, B1 => 
                           data_in(39), B2 => n9_port, Y => n103);
   U111 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_40_port, A2 => n3, B1 => 
                           data_in(40), B2 => n7_port, Y => n101);
   U112 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_41_port, A2 => n3, B1 => 
                           data_in(41), B2 => n7_port, Y => n99);
   U113 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_42_port, A2 => n3, B1 => 
                           data_in(42), B2 => n7_port, Y => n97);
   U114 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_43_port, A2 => n3, B1 => 
                           data_in(43), B2 => n7_port, Y => n95);
   U115 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_44_port, A2 => n3, B1 => 
                           data_in(44), B2 => n7_port, Y => n93);
   U116 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_45_port, A2 => n3, B1 => 
                           data_in(45), B2 => n7_port, Y => n91);
   U117 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_46_port, A2 => n3, B1 => 
                           data_in(46), B2 => n7_port, Y => n89);
   U118 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_47_port, A2 => n3, B1 => 
                           data_in(47), B2 => n7_port, Y => n87);
   U119 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_48_port, A2 => n3, B1 => 
                           data_in(48), B2 => n7_port, Y => n85);
   U120 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_49_port, A2 => n3, B1 => 
                           data_in(49), B2 => n7_port, Y => n83);
   U121 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_50_port, A2 => n3, B1 => 
                           data_in(50), B2 => n7_port, Y => n81);
   U122 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_51_port, A2 => n3, B1 => 
                           data_in(51), B2 => n7_port, Y => n79);
   U123 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_52_port, A2 => n3, B1 => 
                           data_in(52), B2 => n5, Y => n77);
   U124 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_53_port, A2 => n3, B1 => 
                           data_in(53), B2 => n5, Y => n75);
   U125 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_54_port, A2 => n3, B1 => 
                           data_in(54), B2 => n5, Y => n73);
   U126 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_55_port, A2 => n3, B1 => 
                           data_in(55), B2 => n5, Y => n71);
   U127 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_56_port, A2 => n3, B1 => 
                           data_in(56), B2 => n5, Y => n69);
   U128 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_57_port, A2 => n3, B1 => 
                           data_in(57), B2 => n5, Y => n67);
   U129 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_58_port, A2 => n3, B1 => 
                           data_in(58), B2 => n5, Y => n65);
   U130 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_59_port, A2 => n3, B1 => 
                           data_in(59), B2 => n5, Y => n63);
   U131 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_60_port, A2 => n3, B1 => 
                           data_in(60), B2 => n5, Y => n61);
   U132 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_61_port, A2 => n3, B1 => 
                           data_in(61), B2 => n5, Y => n59);
   U133 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_62_port, A2 => n3, B1 => 
                           data_in(62), B2 => n5, Y => n57);
   U134 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_63_port, A2 => n3, B1 => 
                           data_in(63), B2 => n5, Y => n55);
   U136 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N7, Y => n236);
   U137 : OAI22xp5_ASAP7_75t_R port map( A1 => n31, A2 => read_en, B1 => n43, 
                           B2 => n45, Y => n53);
   U139 : OAI22xp5_ASAP7_75t_R port map( A1 => N9, A2 => n49, B1 => write_en, 
                           B2 => N7, Y => n51);
   write_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK 
                           => clk, RESET => n47, SET => n1, QN => N7);
   fifo_reg_1_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n55, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_63_port);
   fifo_reg_1_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n57, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_62_port);
   fifo_reg_1_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n59, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_61_port);
   fifo_reg_1_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n61, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_60_port);
   fifo_reg_0_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n171, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_63_port);
   fifo_reg_0_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n172, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_62_port);
   fifo_reg_0_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n173, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_61_port);
   fifo_reg_0_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n174, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_60_port);
   fifo_reg_1_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n167, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_3_port);
   fifo_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n168, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_2_port);
   fifo_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n169, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_1_port);
   fifo_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n170, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_0_port);
   fifo_reg_1_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n63, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_59_port);
   fifo_reg_1_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n65, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_58_port);
   fifo_reg_1_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n67, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_57_port);
   fifo_reg_1_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n69, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_56_port);
   fifo_reg_1_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n71, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_55_port);
   fifo_reg_1_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n73, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_54_port);
   fifo_reg_1_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n75, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_53_port);
   fifo_reg_1_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n77, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_52_port);
   fifo_reg_1_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_51_port);
   fifo_reg_1_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_50_port);
   fifo_reg_1_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_49_port);
   fifo_reg_1_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_48_port);
   fifo_reg_1_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_47_port);
   fifo_reg_1_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_46_port);
   fifo_reg_1_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_45_port);
   fifo_reg_1_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_44_port);
   fifo_reg_1_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_43_port);
   fifo_reg_1_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_42_port);
   fifo_reg_1_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_41_port);
   fifo_reg_1_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_40_port);
   fifo_reg_1_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_39_port);
   fifo_reg_1_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_38_port);
   fifo_reg_1_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_37_port);
   fifo_reg_1_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_36_port);
   fifo_reg_1_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_35_port);
   fifo_reg_1_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_34_port);
   fifo_reg_1_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n115, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_33_port);
   fifo_reg_1_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n117, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_32_port);
   fifo_reg_1_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n119, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_31_port);
   fifo_reg_1_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n121, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_30_port);
   fifo_reg_1_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n123, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_29_port);
   fifo_reg_1_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n125, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_28_port);
   fifo_reg_1_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n127, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_27_port);
   fifo_reg_1_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n129, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_26_port);
   fifo_reg_1_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n131, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_25_port);
   fifo_reg_1_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n133, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_24_port);
   fifo_reg_1_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n135, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_23_port);
   fifo_reg_1_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n137, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_22_port);
   fifo_reg_1_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n139, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_21_port);
   fifo_reg_1_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n141, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_20_port);
   fifo_reg_1_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n143, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_19_port);
   fifo_reg_1_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n145, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_18_port);
   fifo_reg_1_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n147, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_17_port);
   fifo_reg_1_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n149, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_16_port);
   fifo_reg_1_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n151, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_15_port);
   fifo_reg_1_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n153, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_14_port);
   fifo_reg_1_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n155, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_13_port);
   fifo_reg_1_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n157, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_12_port);
   fifo_reg_1_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n159, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_11_port);
   fifo_reg_1_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n160, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_10_port);
   fifo_reg_1_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n161, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_9_port);
   fifo_reg_1_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n162, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_8_port);
   fifo_reg_1_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n163, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_7_port);
   fifo_reg_1_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n164, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_6_port);
   fifo_reg_1_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n165, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_5_port);
   fifo_reg_1_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n166, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_4_port);
   fifo_reg_0_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n231, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_3_port);
   fifo_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n232, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_2_port);
   fifo_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n233, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_1_port);
   fifo_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n234, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_0_port);
   fifo_reg_0_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n175, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_59_port);
   fifo_reg_0_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n176, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_58_port);
   fifo_reg_0_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n177, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_57_port);
   fifo_reg_0_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n178, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_56_port);
   fifo_reg_0_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n179, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_55_port);
   fifo_reg_0_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n180, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_54_port);
   fifo_reg_0_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n181, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_53_port);
   fifo_reg_0_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n182, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_52_port);
   fifo_reg_0_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n183, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_51_port);
   fifo_reg_0_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n184, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_50_port);
   fifo_reg_0_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n185, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_49_port);
   fifo_reg_0_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n186, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_48_port);
   fifo_reg_0_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n187, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_47_port);
   fifo_reg_0_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n188, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_46_port);
   fifo_reg_0_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n189, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_45_port);
   fifo_reg_0_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n190, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_44_port);
   fifo_reg_0_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n191, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_43_port);
   fifo_reg_0_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n192, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_42_port);
   fifo_reg_0_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n193, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_41_port);
   fifo_reg_0_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n194, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_40_port);
   fifo_reg_0_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n195, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_39_port);
   fifo_reg_0_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n196, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_38_port);
   fifo_reg_0_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n197, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_37_port);
   fifo_reg_0_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n198, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_36_port);
   fifo_reg_0_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n199, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_35_port);
   fifo_reg_0_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n200, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_34_port);
   fifo_reg_0_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n201, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_33_port);
   fifo_reg_0_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n202, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_32_port);
   fifo_reg_0_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n203, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_31_port);
   fifo_reg_0_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n204, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_30_port);
   fifo_reg_0_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n205, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_29_port);
   fifo_reg_0_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n206, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_28_port);
   fifo_reg_0_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n207, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_27_port);
   fifo_reg_0_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n208, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_26_port);
   fifo_reg_0_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n209, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_25_port);
   fifo_reg_0_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n210, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_24_port);
   fifo_reg_0_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n211, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_23_port);
   fifo_reg_0_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n212, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_22_port);
   fifo_reg_0_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n213, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_21_port);
   fifo_reg_0_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n214, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_20_port);
   fifo_reg_0_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n215, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_19_port);
   fifo_reg_0_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n216, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_18_port);
   fifo_reg_0_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n217, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_17_port);
   fifo_reg_0_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n218, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_16_port);
   fifo_reg_0_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n219, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_15_port);
   fifo_reg_0_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n220, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_14_port);
   fifo_reg_0_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n221, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_13_port);
   fifo_reg_0_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n222, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_12_port);
   fifo_reg_0_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n223, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_11_port);
   fifo_reg_0_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n224, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_10_port);
   fifo_reg_0_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n225, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_9_port);
   fifo_reg_0_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n226, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_8_port);
   fifo_reg_0_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n227, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_7_port);
   fifo_reg_0_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n228, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_6_port);
   fifo_reg_0_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n229, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_5_port);
   fifo_reg_0_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n230, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_4_port);
   valid_data_reg : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n235, CLK => clk, 
                           RESET => n47, SET => n1, QN => valid_data_port);
   read_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK 
                           => clk, RESET => n47, SET => n1, QN => 
                           read_pointer_0_port);
   U69 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U135 : INVx3_ASAP7_75t_R port map( A => rst, Y => n47);
   U138 : INVx1_ASAP7_75t_R port map( A => read_en, Y => n45);
   U140 : INVx1_ASAP7_75t_R port map( A => n29, Y => n17);
   U141 : INVx1_ASAP7_75t_R port map( A => n15, Y => n3);
   U142 : INVx1_ASAP7_75t_R port map( A => n31, Y => n43);
   U207 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n29);
   U208 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n15);
   U209 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n27);
   U210 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n25);
   U211 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n23);
   U212 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n21);
   U213 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n19);
   U214 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n13);
   U215 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n11);
   U216 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n9_port);
   U217 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n7_port);
   U218 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n5);
   U219 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n31);
   U220 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n33);
   U221 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n41);
   U222 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n39);
   U223 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n37);
   U224 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n35);
   U225 : INVx1_ASAP7_75t_R port map( A => N7, Y => N9);
   U226 : INVx1_ASAP7_75t_R port map( A => write_en, Y => n49);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity fifo_buff_depth2_6 is

   port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, clk, 
         rst : in std_logic;  data_out : out std_logic_vector (63 downto 0);  
         valid_data : out std_logic);

end fifo_buff_depth2_6;

architecture SYN_rtl of fifo_buff_depth2_6 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx3_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal valid_data_port, read_pointer_0_port, fifo_1_63_port, fifo_1_62_port,
      fifo_1_61_port, fifo_1_60_port, fifo_1_59_port, fifo_1_58_port, 
      fifo_1_57_port, fifo_1_56_port, fifo_1_55_port, fifo_1_54_port, 
      fifo_1_53_port, fifo_1_52_port, fifo_1_51_port, fifo_1_50_port, 
      fifo_1_49_port, fifo_1_48_port, fifo_1_47_port, fifo_1_46_port, 
      fifo_1_45_port, fifo_1_44_port, fifo_1_43_port, fifo_1_42_port, 
      fifo_1_41_port, fifo_1_40_port, fifo_1_39_port, fifo_1_38_port, 
      fifo_1_37_port, fifo_1_36_port, fifo_1_35_port, fifo_1_34_port, 
      fifo_1_33_port, fifo_1_32_port, fifo_1_31_port, fifo_1_30_port, 
      fifo_1_29_port, fifo_1_28_port, fifo_1_27_port, fifo_1_26_port, 
      fifo_1_25_port, fifo_1_24_port, fifo_1_23_port, fifo_1_22_port, 
      fifo_1_21_port, fifo_1_20_port, fifo_1_19_port, fifo_1_18_port, 
      fifo_1_17_port, fifo_1_16_port, fifo_1_15_port, fifo_1_14_port, 
      fifo_1_13_port, fifo_1_12_port, fifo_1_11_port, fifo_1_10_port, 
      fifo_1_9_port, fifo_1_8_port, fifo_1_7_port, fifo_1_6_port, fifo_1_5_port
      , fifo_1_4_port, fifo_1_3_port, fifo_1_2_port, fifo_1_1_port, 
      fifo_1_0_port, fifo_0_63_port, fifo_0_62_port, fifo_0_61_port, 
      fifo_0_60_port, fifo_0_59_port, fifo_0_58_port, fifo_0_57_port, 
      fifo_0_56_port, fifo_0_55_port, fifo_0_54_port, fifo_0_53_port, 
      fifo_0_52_port, fifo_0_51_port, fifo_0_50_port, fifo_0_49_port, 
      fifo_0_48_port, fifo_0_47_port, fifo_0_46_port, fifo_0_45_port, 
      fifo_0_44_port, fifo_0_43_port, fifo_0_42_port, fifo_0_41_port, 
      fifo_0_40_port, fifo_0_39_port, fifo_0_38_port, fifo_0_37_port, 
      fifo_0_36_port, fifo_0_35_port, fifo_0_34_port, fifo_0_33_port, 
      fifo_0_32_port, fifo_0_31_port, fifo_0_30_port, fifo_0_29_port, 
      fifo_0_28_port, fifo_0_27_port, fifo_0_26_port, fifo_0_25_port, 
      fifo_0_24_port, fifo_0_23_port, fifo_0_22_port, fifo_0_21_port, 
      fifo_0_20_port, fifo_0_19_port, fifo_0_18_port, fifo_0_17_port, 
      fifo_0_16_port, fifo_0_15_port, fifo_0_14_port, fifo_0_13_port, 
      fifo_0_12_port, fifo_0_11_port, fifo_0_10_port, fifo_0_9_port, 
      fifo_0_8_port, fifo_0_7_port, fifo_0_6_port, fifo_0_5_port, fifo_0_4_port
      , fifo_0_3_port, fifo_0_2_port, fifo_0_1_port, fifo_0_0_port, N7, N9, n1,
      n3, n5, n7_port, n9_port, n11, n13, n15, n17, n19, n21, n23, n25, n27, 
      n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57
      , n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, 
      n87, n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, n111, 
      n113, n115, n117, n119, n121, n123, n125, n127, n129, n131, n133, n135, 
      n137, n139, n141, n143, n145, n147, n149, n151, n153, n155, n157, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238 : std_logic;

begin
   valid_data <= valid_data_port;
   
   U4 : XOR2xp5_ASAP7_75t_R port map( A => N7, B => n43, Y => n238);
   U143 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_9_port, B1 => 
                           n43, B2 => fifo_0_9_port, Y => data_out(9));
   U144 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_8_port, B1 => 
                           n43, B2 => fifo_0_8_port, Y => data_out(8));
   U145 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_7_port, B1 => 
                           n43, B2 => fifo_0_7_port, Y => data_out(7));
   U146 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_6_port, B1 => 
                           n43, B2 => fifo_0_6_port, Y => data_out(6));
   U147 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_63_port, B1 => 
                           n43, B2 => fifo_0_63_port, Y => data_out(63));
   U148 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_62_port, B1 => 
                           n43, B2 => fifo_0_62_port, Y => data_out(62));
   U149 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_61_port, B1 => 
                           n43, B2 => fifo_0_61_port, Y => data_out(61));
   U150 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_60_port, B1 => 
                           n43, B2 => fifo_0_60_port, Y => data_out(60));
   U151 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_5_port, B1 => 
                           n43, B2 => fifo_0_5_port, Y => data_out(5));
   U152 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_59_port, B1 => 
                           n43, B2 => fifo_0_59_port, Y => data_out(59));
   U153 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_58_port, B1 => 
                           n43, B2 => fifo_0_58_port, Y => data_out(58));
   U154 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_57_port, B1 => 
                           n43, B2 => fifo_0_57_port, Y => data_out(57));
   U155 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_56_port, B1 => 
                           n43, B2 => fifo_0_56_port, Y => data_out(56));
   U156 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_55_port, B1 => 
                           n43, B2 => fifo_0_55_port, Y => data_out(55));
   U157 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_54_port, B1 => 
                           n43, B2 => fifo_0_54_port, Y => data_out(54));
   U158 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_53_port, B1 => 
                           n43, B2 => fifo_0_53_port, Y => data_out(53));
   U159 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_52_port, B1 => 
                           n43, B2 => fifo_0_52_port, Y => data_out(52));
   U160 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_51_port, B1 => 
                           n43, B2 => fifo_0_51_port, Y => data_out(51));
   U161 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_50_port, B1 => 
                           n43, B2 => fifo_0_50_port, Y => data_out(50));
   U162 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_4_port, B1 => 
                           n43, B2 => fifo_0_4_port, Y => data_out(4));
   U163 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_49_port, B1 => 
                           n43, B2 => fifo_0_49_port, Y => data_out(49));
   U164 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_48_port, B1 => 
                           n43, B2 => fifo_0_48_port, Y => data_out(48));
   U165 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_47_port, B1 => 
                           n43, B2 => fifo_0_47_port, Y => data_out(47));
   U166 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_46_port, B1 => 
                           n43, B2 => fifo_0_46_port, Y => data_out(46));
   U167 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_45_port, B1 => 
                           n43, B2 => fifo_0_45_port, Y => data_out(45));
   U168 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_44_port, B1 => 
                           n43, B2 => fifo_0_44_port, Y => data_out(44));
   U169 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_43_port, B1 => 
                           n43, B2 => fifo_0_43_port, Y => data_out(43));
   U170 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_42_port, B1 => 
                           n43, B2 => fifo_0_42_port, Y => data_out(42));
   U171 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_41_port, B1 => 
                           n43, B2 => fifo_0_41_port, Y => data_out(41));
   U172 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_40_port, B1 => 
                           n43, B2 => fifo_0_40_port, Y => data_out(40));
   U173 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_3_port, B1 => 
                           n43, B2 => fifo_0_3_port, Y => data_out(3));
   U174 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_39_port, B1 => 
                           n43, B2 => fifo_0_39_port, Y => data_out(39));
   U175 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_38_port, B1 => 
                           n43, B2 => fifo_0_38_port, Y => data_out(38));
   U176 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_37_port, B1 => 
                           n43, B2 => fifo_0_37_port, Y => data_out(37));
   U177 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_36_port, B1 => 
                           n43, B2 => fifo_0_36_port, Y => data_out(36));
   U178 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_35_port, B1 => 
                           n43, B2 => fifo_0_35_port, Y => data_out(35));
   U179 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_34_port, B1 => 
                           n43, B2 => fifo_0_34_port, Y => data_out(34));
   U180 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_33_port, B1 => 
                           n43, B2 => fifo_0_33_port, Y => data_out(33));
   U181 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_32_port, B1 => 
                           n43, B2 => fifo_0_32_port, Y => data_out(32));
   U182 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_31_port, B1 => 
                           n43, B2 => fifo_0_31_port, Y => data_out(31));
   U183 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_30_port, B1 => 
                           n43, B2 => fifo_0_30_port, Y => data_out(30));
   U184 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_2_port, B1 => 
                           n43, B2 => fifo_0_2_port, Y => data_out(2));
   U185 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_29_port, B1 => 
                           n43, B2 => fifo_0_29_port, Y => data_out(29));
   U186 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_28_port, B1 => 
                           n43, B2 => fifo_0_28_port, Y => data_out(28));
   U187 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_27_port, B1 => 
                           n43, B2 => fifo_0_27_port, Y => data_out(27));
   U188 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_26_port, B1 => 
                           n43, B2 => fifo_0_26_port, Y => data_out(26));
   U189 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_25_port, B1 => 
                           n43, B2 => fifo_0_25_port, Y => data_out(25));
   U190 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_24_port, B1 => 
                           n43, B2 => fifo_0_24_port, Y => data_out(24));
   U191 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_23_port, B1 => 
                           n43, B2 => fifo_0_23_port, Y => data_out(23));
   U192 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_22_port, B1 => 
                           n43, B2 => fifo_0_22_port, Y => data_out(22));
   U193 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_21_port, B1 => 
                           n43, B2 => fifo_0_21_port, Y => data_out(21));
   U194 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_20_port, B1 => 
                           n43, B2 => fifo_0_20_port, Y => data_out(20));
   U195 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_1_port, B1 => 
                           n43, B2 => fifo_0_1_port, Y => data_out(1));
   U196 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_19_port, B1 => 
                           n43, B2 => fifo_0_19_port, Y => data_out(19));
   U197 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_18_port, B1 => 
                           n43, B2 => fifo_0_18_port, Y => data_out(18));
   U198 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_17_port, B1 => 
                           n43, B2 => fifo_0_17_port, Y => data_out(17));
   U199 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_16_port, B1 => 
                           n43, B2 => fifo_0_16_port, Y => data_out(16));
   U200 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_15_port, B1 => 
                           n43, B2 => fifo_0_15_port, Y => data_out(15));
   U201 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_14_port, B1 => 
                           n43, B2 => fifo_0_14_port, Y => data_out(14));
   U202 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_13_port, B1 => 
                           n43, B2 => fifo_0_13_port, Y => data_out(13));
   U203 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_12_port, B1 => 
                           n43, B2 => fifo_0_12_port, Y => data_out(12));
   U204 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_11_port, B1 => 
                           n43, B2 => fifo_0_11_port, Y => data_out(11));
   U205 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_10_port, B1 => 
                           n43, B2 => fifo_0_10_port, Y => data_out(10));
   U206 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_0_port, B1 => 
                           n43, B2 => fifo_0_0_port, Y => data_out(0));
   U3 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n47, A2 => n238, B => 
                           valid_data_port, C => write_en, Y => n235);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_0_port, A2 => n17, B1 => 
                           data_in(0), B2 => n29, Y => n234);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_1_port, A2 => n17, B1 => 
                           data_in(1), B2 => n29, Y => n233);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_2_port, A2 => n17, B1 => 
                           data_in(2), B2 => n29, Y => n232);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_3_port, A2 => n17, B1 => 
                           data_in(3), B2 => n29, Y => n231);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_4_port, A2 => n17, B1 => 
                           data_in(4), B2 => n27, Y => n230);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_5_port, A2 => n17, B1 => 
                           data_in(5), B2 => n27, Y => n229);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_6_port, A2 => n17, B1 => 
                           data_in(6), B2 => n27, Y => n228);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_7_port, A2 => n17, B1 => 
                           data_in(7), B2 => n27, Y => n227);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_8_port, A2 => n17, B1 => 
                           data_in(8), B2 => n27, Y => n226);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_9_port, A2 => n17, B1 => 
                           data_in(9), B2 => n27, Y => n225);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_10_port, A2 => n17, B1 => 
                           data_in(10), B2 => n27, Y => n224);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_11_port, A2 => n17, B1 => 
                           data_in(11), B2 => n27, Y => n223);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_12_port, A2 => n17, B1 => 
                           data_in(12), B2 => n27, Y => n222);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_13_port, A2 => n17, B1 => 
                           data_in(13), B2 => n27, Y => n221);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_14_port, A2 => n17, B1 => 
                           data_in(14), B2 => n27, Y => n220);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_15_port, A2 => n17, B1 => 
                           data_in(15), B2 => n27, Y => n219);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_16_port, A2 => n17, B1 => 
                           data_in(16), B2 => n25, Y => n218);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_17_port, A2 => n17, B1 => 
                           data_in(17), B2 => n25, Y => n217);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_18_port, A2 => n17, B1 => 
                           data_in(18), B2 => n25, Y => n216);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_19_port, A2 => n17, B1 => 
                           data_in(19), B2 => n25, Y => n215);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_20_port, A2 => n17, B1 => 
                           data_in(20), B2 => n25, Y => n214);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_21_port, A2 => n17, B1 => 
                           data_in(21), B2 => n25, Y => n213);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_22_port, A2 => n17, B1 => 
                           data_in(22), B2 => n25, Y => n212);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_23_port, A2 => n17, B1 => 
                           data_in(23), B2 => n25, Y => n211);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_24_port, A2 => n17, B1 => 
                           data_in(24), B2 => n25, Y => n210);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_25_port, A2 => n17, B1 => 
                           data_in(25), B2 => n25, Y => n209);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_26_port, A2 => n17, B1 => 
                           data_in(26), B2 => n25, Y => n208);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_27_port, A2 => n17, B1 => 
                           data_in(27), B2 => n25, Y => n207);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_28_port, A2 => n17, B1 => 
                           data_in(28), B2 => n23, Y => n206);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_29_port, A2 => n17, B1 => 
                           data_in(29), B2 => n23, Y => n205);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_30_port, A2 => n17, B1 => 
                           data_in(30), B2 => n23, Y => n204);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_31_port, A2 => n17, B1 => 
                           data_in(31), B2 => n23, Y => n203);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_32_port, A2 => n17, B1 => 
                           data_in(32), B2 => n23, Y => n202);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_33_port, A2 => n17, B1 => 
                           data_in(33), B2 => n23, Y => n201);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_34_port, A2 => n17, B1 => 
                           data_in(34), B2 => n23, Y => n200);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_35_port, A2 => n17, B1 => 
                           data_in(35), B2 => n23, Y => n199);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_36_port, A2 => n17, B1 => 
                           data_in(36), B2 => n23, Y => n198);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_37_port, A2 => n17, B1 => 
                           data_in(37), B2 => n23, Y => n197);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_38_port, A2 => n17, B1 => 
                           data_in(38), B2 => n23, Y => n196);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_39_port, A2 => n17, B1 => 
                           data_in(39), B2 => n23, Y => n195);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_40_port, A2 => n17, B1 => 
                           data_in(40), B2 => n21, Y => n194);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_41_port, A2 => n17, B1 => 
                           data_in(41), B2 => n21, Y => n193);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_42_port, A2 => n17, B1 => 
                           data_in(42), B2 => n21, Y => n192);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_43_port, A2 => n17, B1 => 
                           data_in(43), B2 => n21, Y => n191);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_44_port, A2 => n17, B1 => 
                           data_in(44), B2 => n21, Y => n190);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_45_port, A2 => n17, B1 => 
                           data_in(45), B2 => n21, Y => n189);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_46_port, A2 => n17, B1 => 
                           data_in(46), B2 => n21, Y => n188);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_47_port, A2 => n17, B1 => 
                           data_in(47), B2 => n21, Y => n187);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_48_port, A2 => n17, B1 => 
                           data_in(48), B2 => n21, Y => n186);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_49_port, A2 => n17, B1 => 
                           data_in(49), B2 => n21, Y => n185);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_50_port, A2 => n17, B1 => 
                           data_in(50), B2 => n21, Y => n184);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_51_port, A2 => n17, B1 => 
                           data_in(51), B2 => n21, Y => n183);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_52_port, A2 => n17, B1 => 
                           data_in(52), B2 => n19, Y => n182);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_53_port, A2 => n17, B1 => 
                           data_in(53), B2 => n19, Y => n181);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_54_port, A2 => n17, B1 => 
                           data_in(54), B2 => n19, Y => n180);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_55_port, A2 => n17, B1 => 
                           data_in(55), B2 => n19, Y => n179);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_56_port, A2 => n17, B1 => 
                           data_in(56), B2 => n19, Y => n178);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_57_port, A2 => n17, B1 => 
                           data_in(57), B2 => n19, Y => n177);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_58_port, A2 => n17, B1 => 
                           data_in(58), B2 => n19, Y => n176);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_59_port, A2 => n17, B1 => 
                           data_in(59), B2 => n19, Y => n175);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_60_port, A2 => n17, B1 => 
                           data_in(60), B2 => n19, Y => n174);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_61_port, A2 => n17, B1 => 
                           data_in(61), B2 => n19, Y => n173);
   U67 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_62_port, A2 => n17, B1 => 
                           data_in(62), B2 => n19, Y => n172);
   U68 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_63_port, A2 => n17, B1 => 
                           data_in(63), B2 => n19, Y => n171);
   U70 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N9, Y => n237);
   U71 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_0_port, A2 => n3, B1 => 
                           data_in(0), B2 => n15, Y => n170);
   U72 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_1_port, A2 => n3, B1 => 
                           data_in(1), B2 => n15, Y => n169);
   U73 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_2_port, A2 => n3, B1 => 
                           data_in(2), B2 => n15, Y => n168);
   U74 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_3_port, A2 => n3, B1 => 
                           data_in(3), B2 => n15, Y => n167);
   U75 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_4_port, A2 => n3, B1 => 
                           data_in(4), B2 => n13, Y => n166);
   U76 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_5_port, A2 => n3, B1 => 
                           data_in(5), B2 => n13, Y => n165);
   U77 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_6_port, A2 => n3, B1 => 
                           data_in(6), B2 => n13, Y => n164);
   U78 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_7_port, A2 => n3, B1 => 
                           data_in(7), B2 => n13, Y => n163);
   U79 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_8_port, A2 => n3, B1 => 
                           data_in(8), B2 => n13, Y => n162);
   U80 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_9_port, A2 => n3, B1 => 
                           data_in(9), B2 => n13, Y => n161);
   U81 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_10_port, A2 => n3, B1 => 
                           data_in(10), B2 => n13, Y => n160);
   U82 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_11_port, A2 => n3, B1 => 
                           data_in(11), B2 => n13, Y => n159);
   U83 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_12_port, A2 => n3, B1 => 
                           data_in(12), B2 => n13, Y => n157);
   U84 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_13_port, A2 => n3, B1 => 
                           data_in(13), B2 => n13, Y => n155);
   U85 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_14_port, A2 => n3, B1 => 
                           data_in(14), B2 => n13, Y => n153);
   U86 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_15_port, A2 => n3, B1 => 
                           data_in(15), B2 => n13, Y => n151);
   U87 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_16_port, A2 => n3, B1 => 
                           data_in(16), B2 => n11, Y => n149);
   U88 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_17_port, A2 => n3, B1 => 
                           data_in(17), B2 => n11, Y => n147);
   U89 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_18_port, A2 => n3, B1 => 
                           data_in(18), B2 => n11, Y => n145);
   U90 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_19_port, A2 => n3, B1 => 
                           data_in(19), B2 => n11, Y => n143);
   U91 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_20_port, A2 => n3, B1 => 
                           data_in(20), B2 => n11, Y => n141);
   U92 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_21_port, A2 => n3, B1 => 
                           data_in(21), B2 => n11, Y => n139);
   U93 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_22_port, A2 => n3, B1 => 
                           data_in(22), B2 => n11, Y => n137);
   U94 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_23_port, A2 => n3, B1 => 
                           data_in(23), B2 => n11, Y => n135);
   U95 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_24_port, A2 => n3, B1 => 
                           data_in(24), B2 => n11, Y => n133);
   U96 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_25_port, A2 => n3, B1 => 
                           data_in(25), B2 => n11, Y => n131);
   U97 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_26_port, A2 => n3, B1 => 
                           data_in(26), B2 => n11, Y => n129);
   U98 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_27_port, A2 => n3, B1 => 
                           data_in(27), B2 => n11, Y => n127);
   U99 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_28_port, A2 => n3, B1 => 
                           data_in(28), B2 => n9_port, Y => n125);
   U100 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_29_port, A2 => n3, B1 => 
                           data_in(29), B2 => n9_port, Y => n123);
   U101 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_30_port, A2 => n3, B1 => 
                           data_in(30), B2 => n9_port, Y => n121);
   U102 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_31_port, A2 => n3, B1 => 
                           data_in(31), B2 => n9_port, Y => n119);
   U103 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_32_port, A2 => n3, B1 => 
                           data_in(32), B2 => n9_port, Y => n117);
   U104 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_33_port, A2 => n3, B1 => 
                           data_in(33), B2 => n9_port, Y => n115);
   U105 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_34_port, A2 => n3, B1 => 
                           data_in(34), B2 => n9_port, Y => n113);
   U106 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_35_port, A2 => n3, B1 => 
                           data_in(35), B2 => n9_port, Y => n111);
   U107 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_36_port, A2 => n3, B1 => 
                           data_in(36), B2 => n9_port, Y => n109);
   U108 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_37_port, A2 => n3, B1 => 
                           data_in(37), B2 => n9_port, Y => n107);
   U109 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_38_port, A2 => n3, B1 => 
                           data_in(38), B2 => n9_port, Y => n105);
   U110 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_39_port, A2 => n3, B1 => 
                           data_in(39), B2 => n9_port, Y => n103);
   U111 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_40_port, A2 => n3, B1 => 
                           data_in(40), B2 => n7_port, Y => n101);
   U112 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_41_port, A2 => n3, B1 => 
                           data_in(41), B2 => n7_port, Y => n99);
   U113 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_42_port, A2 => n3, B1 => 
                           data_in(42), B2 => n7_port, Y => n97);
   U114 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_43_port, A2 => n3, B1 => 
                           data_in(43), B2 => n7_port, Y => n95);
   U115 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_44_port, A2 => n3, B1 => 
                           data_in(44), B2 => n7_port, Y => n93);
   U116 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_45_port, A2 => n3, B1 => 
                           data_in(45), B2 => n7_port, Y => n91);
   U117 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_46_port, A2 => n3, B1 => 
                           data_in(46), B2 => n7_port, Y => n89);
   U118 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_47_port, A2 => n3, B1 => 
                           data_in(47), B2 => n7_port, Y => n87);
   U119 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_48_port, A2 => n3, B1 => 
                           data_in(48), B2 => n7_port, Y => n85);
   U120 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_49_port, A2 => n3, B1 => 
                           data_in(49), B2 => n7_port, Y => n83);
   U121 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_50_port, A2 => n3, B1 => 
                           data_in(50), B2 => n7_port, Y => n81);
   U122 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_51_port, A2 => n3, B1 => 
                           data_in(51), B2 => n7_port, Y => n79);
   U123 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_52_port, A2 => n3, B1 => 
                           data_in(52), B2 => n5, Y => n77);
   U124 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_53_port, A2 => n3, B1 => 
                           data_in(53), B2 => n5, Y => n75);
   U125 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_54_port, A2 => n3, B1 => 
                           data_in(54), B2 => n5, Y => n73);
   U126 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_55_port, A2 => n3, B1 => 
                           data_in(55), B2 => n5, Y => n71);
   U127 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_56_port, A2 => n3, B1 => 
                           data_in(56), B2 => n5, Y => n69);
   U128 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_57_port, A2 => n3, B1 => 
                           data_in(57), B2 => n5, Y => n67);
   U129 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_58_port, A2 => n3, B1 => 
                           data_in(58), B2 => n5, Y => n65);
   U130 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_59_port, A2 => n3, B1 => 
                           data_in(59), B2 => n5, Y => n63);
   U131 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_60_port, A2 => n3, B1 => 
                           data_in(60), B2 => n5, Y => n61);
   U132 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_61_port, A2 => n3, B1 => 
                           data_in(61), B2 => n5, Y => n59);
   U133 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_62_port, A2 => n3, B1 => 
                           data_in(62), B2 => n5, Y => n57);
   U134 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_63_port, A2 => n3, B1 => 
                           data_in(63), B2 => n5, Y => n55);
   U136 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N7, Y => n236);
   U137 : OAI22xp5_ASAP7_75t_R port map( A1 => n31, A2 => read_en, B1 => n43, 
                           B2 => n47, Y => n53);
   U139 : OAI22xp5_ASAP7_75t_R port map( A1 => N9, A2 => n49, B1 => write_en, 
                           B2 => N7, Y => n51);
   write_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK 
                           => clk, RESET => n45, SET => n1, QN => N7);
   fifo_reg_1_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n55, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_63_port);
   fifo_reg_1_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n57, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_62_port);
   fifo_reg_1_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n59, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_61_port);
   fifo_reg_1_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n61, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_60_port);
   fifo_reg_0_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n171, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_63_port);
   fifo_reg_0_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n172, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_62_port);
   fifo_reg_0_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n173, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_61_port);
   fifo_reg_0_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n174, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_60_port);
   fifo_reg_1_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n167, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_3_port);
   fifo_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n168, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_2_port);
   fifo_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n169, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_1_port);
   fifo_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n170, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_0_port);
   fifo_reg_1_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n63, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_59_port);
   fifo_reg_1_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n65, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_58_port);
   fifo_reg_1_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n67, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_57_port);
   fifo_reg_1_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n69, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_56_port);
   fifo_reg_1_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n71, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_55_port);
   fifo_reg_1_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n73, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_54_port);
   fifo_reg_1_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n75, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_53_port);
   fifo_reg_1_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n77, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_52_port);
   fifo_reg_1_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_51_port);
   fifo_reg_1_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_50_port);
   fifo_reg_1_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_49_port);
   fifo_reg_1_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_48_port);
   fifo_reg_1_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_47_port);
   fifo_reg_1_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_46_port);
   fifo_reg_1_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_45_port);
   fifo_reg_1_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_44_port);
   fifo_reg_1_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_43_port);
   fifo_reg_1_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_42_port);
   fifo_reg_1_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_41_port);
   fifo_reg_1_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_40_port);
   fifo_reg_1_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_39_port);
   fifo_reg_1_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_38_port);
   fifo_reg_1_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_37_port);
   fifo_reg_1_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_36_port);
   fifo_reg_1_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_35_port);
   fifo_reg_1_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_34_port);
   fifo_reg_1_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n115, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_33_port);
   fifo_reg_1_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n117, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_32_port);
   fifo_reg_1_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n119, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_31_port);
   fifo_reg_1_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n121, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_30_port);
   fifo_reg_1_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n123, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_29_port);
   fifo_reg_1_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n125, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_28_port);
   fifo_reg_1_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n127, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_27_port);
   fifo_reg_1_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n129, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_26_port);
   fifo_reg_1_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n131, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_25_port);
   fifo_reg_1_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n133, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_24_port);
   fifo_reg_1_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n135, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_23_port);
   fifo_reg_1_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n137, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_22_port);
   fifo_reg_1_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n139, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_21_port);
   fifo_reg_1_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n141, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_20_port);
   fifo_reg_1_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n143, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_19_port);
   fifo_reg_1_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n145, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_18_port);
   fifo_reg_1_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n147, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_17_port);
   fifo_reg_1_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n149, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_16_port);
   fifo_reg_1_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n151, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_15_port);
   fifo_reg_1_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n153, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_14_port);
   fifo_reg_1_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n155, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_13_port);
   fifo_reg_1_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n157, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_12_port);
   fifo_reg_1_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n159, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_11_port);
   fifo_reg_1_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n160, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_10_port);
   fifo_reg_1_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n161, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_9_port);
   fifo_reg_1_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n162, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_8_port);
   fifo_reg_1_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n163, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_7_port);
   fifo_reg_1_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n164, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_6_port);
   fifo_reg_1_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n165, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_5_port);
   fifo_reg_1_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n166, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_4_port);
   fifo_reg_0_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n231, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_3_port);
   fifo_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n232, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_2_port);
   fifo_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n233, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_1_port);
   fifo_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n234, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_0_port);
   fifo_reg_0_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n175, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_59_port);
   fifo_reg_0_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n176, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_58_port);
   fifo_reg_0_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n177, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_57_port);
   fifo_reg_0_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n178, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_56_port);
   fifo_reg_0_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n179, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_55_port);
   fifo_reg_0_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n180, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_54_port);
   fifo_reg_0_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n181, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_53_port);
   fifo_reg_0_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n182, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_52_port);
   fifo_reg_0_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n183, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_51_port);
   fifo_reg_0_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n184, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_50_port);
   fifo_reg_0_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n185, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_49_port);
   fifo_reg_0_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n186, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_48_port);
   fifo_reg_0_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n187, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_47_port);
   fifo_reg_0_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n188, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_46_port);
   fifo_reg_0_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n189, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_45_port);
   fifo_reg_0_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n190, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_44_port);
   fifo_reg_0_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n191, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_43_port);
   fifo_reg_0_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n192, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_42_port);
   fifo_reg_0_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n193, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_41_port);
   fifo_reg_0_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n194, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_40_port);
   fifo_reg_0_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n195, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_39_port);
   fifo_reg_0_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n196, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_38_port);
   fifo_reg_0_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n197, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_37_port);
   fifo_reg_0_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n198, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_36_port);
   fifo_reg_0_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n199, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_35_port);
   fifo_reg_0_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n200, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_34_port);
   fifo_reg_0_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n201, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_33_port);
   fifo_reg_0_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n202, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_32_port);
   fifo_reg_0_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n203, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_31_port);
   fifo_reg_0_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n204, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_30_port);
   fifo_reg_0_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n205, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_29_port);
   fifo_reg_0_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n206, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_28_port);
   fifo_reg_0_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n207, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_27_port);
   fifo_reg_0_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n208, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_26_port);
   fifo_reg_0_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n209, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_25_port);
   fifo_reg_0_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n210, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_24_port);
   fifo_reg_0_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n211, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_23_port);
   fifo_reg_0_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n212, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_22_port);
   fifo_reg_0_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n213, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_21_port);
   fifo_reg_0_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n214, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_20_port);
   fifo_reg_0_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n215, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_19_port);
   fifo_reg_0_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n216, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_18_port);
   fifo_reg_0_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n217, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_17_port);
   fifo_reg_0_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n218, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_16_port);
   fifo_reg_0_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n219, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_15_port);
   fifo_reg_0_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n220, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_14_port);
   fifo_reg_0_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n221, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_13_port);
   fifo_reg_0_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n222, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_12_port);
   fifo_reg_0_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n223, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_11_port);
   fifo_reg_0_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n224, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_10_port);
   fifo_reg_0_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n225, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_9_port);
   fifo_reg_0_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n226, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_8_port);
   fifo_reg_0_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n227, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_7_port);
   fifo_reg_0_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n228, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_6_port);
   fifo_reg_0_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n229, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_5_port);
   fifo_reg_0_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n230, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_4_port);
   read_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK 
                           => clk, RESET => n45, SET => n1, QN => 
                           read_pointer_0_port);
   valid_data_reg : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n235, CLK => clk, 
                           RESET => n45, SET => n1, QN => valid_data_port);
   U69 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U135 : INVx3_ASAP7_75t_R port map( A => rst, Y => n45);
   U138 : INVx1_ASAP7_75t_R port map( A => n29, Y => n17);
   U140 : INVx1_ASAP7_75t_R port map( A => n15, Y => n3);
   U141 : INVx1_ASAP7_75t_R port map( A => n31, Y => n43);
   U142 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n29);
   U207 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n15);
   U208 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n27);
   U209 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n25);
   U210 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n23);
   U211 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n21);
   U212 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n19);
   U213 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n13);
   U214 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n11);
   U215 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n9_port);
   U216 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n7_port);
   U217 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n5);
   U218 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n31);
   U219 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n33);
   U220 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n41);
   U221 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n39);
   U222 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n37);
   U223 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n35);
   U224 : INVx1_ASAP7_75t_R port map( A => read_en, Y => n47);
   U225 : INVx1_ASAP7_75t_R port map( A => N7, Y => N9);
   U226 : INVx1_ASAP7_75t_R port map( A => write_en, Y => n49);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity fifo_buff_depth2_5 is

   port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, clk, 
         rst : in std_logic;  data_out : out std_logic_vector (63 downto 0);  
         valid_data : out std_logic);

end fifo_buff_depth2_5;

architecture SYN_rtl of fifo_buff_depth2_5 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx3_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal valid_data_port, read_pointer_0_port, fifo_1_63_port, fifo_1_62_port,
      fifo_1_61_port, fifo_1_60_port, fifo_1_59_port, fifo_1_58_port, 
      fifo_1_57_port, fifo_1_56_port, fifo_1_55_port, fifo_1_54_port, 
      fifo_1_53_port, fifo_1_52_port, fifo_1_51_port, fifo_1_50_port, 
      fifo_1_49_port, fifo_1_48_port, fifo_1_47_port, fifo_1_46_port, 
      fifo_1_45_port, fifo_1_44_port, fifo_1_43_port, fifo_1_42_port, 
      fifo_1_41_port, fifo_1_40_port, fifo_1_39_port, fifo_1_38_port, 
      fifo_1_37_port, fifo_1_36_port, fifo_1_35_port, fifo_1_34_port, 
      fifo_1_33_port, fifo_1_32_port, fifo_1_31_port, fifo_1_30_port, 
      fifo_1_29_port, fifo_1_28_port, fifo_1_27_port, fifo_1_26_port, 
      fifo_1_25_port, fifo_1_24_port, fifo_1_23_port, fifo_1_22_port, 
      fifo_1_21_port, fifo_1_20_port, fifo_1_19_port, fifo_1_18_port, 
      fifo_1_17_port, fifo_1_16_port, fifo_1_15_port, fifo_1_14_port, 
      fifo_1_13_port, fifo_1_12_port, fifo_1_11_port, fifo_1_10_port, 
      fifo_1_9_port, fifo_1_8_port, fifo_1_7_port, fifo_1_6_port, fifo_1_5_port
      , fifo_1_4_port, fifo_1_3_port, fifo_1_2_port, fifo_1_1_port, 
      fifo_1_0_port, fifo_0_63_port, fifo_0_62_port, fifo_0_61_port, 
      fifo_0_60_port, fifo_0_59_port, fifo_0_58_port, fifo_0_57_port, 
      fifo_0_56_port, fifo_0_55_port, fifo_0_54_port, fifo_0_53_port, 
      fifo_0_52_port, fifo_0_51_port, fifo_0_50_port, fifo_0_49_port, 
      fifo_0_48_port, fifo_0_47_port, fifo_0_46_port, fifo_0_45_port, 
      fifo_0_44_port, fifo_0_43_port, fifo_0_42_port, fifo_0_41_port, 
      fifo_0_40_port, fifo_0_39_port, fifo_0_38_port, fifo_0_37_port, 
      fifo_0_36_port, fifo_0_35_port, fifo_0_34_port, fifo_0_33_port, 
      fifo_0_32_port, fifo_0_31_port, fifo_0_30_port, fifo_0_29_port, 
      fifo_0_28_port, fifo_0_27_port, fifo_0_26_port, fifo_0_25_port, 
      fifo_0_24_port, fifo_0_23_port, fifo_0_22_port, fifo_0_21_port, 
      fifo_0_20_port, fifo_0_19_port, fifo_0_18_port, fifo_0_17_port, 
      fifo_0_16_port, fifo_0_15_port, fifo_0_14_port, fifo_0_13_port, 
      fifo_0_12_port, fifo_0_11_port, fifo_0_10_port, fifo_0_9_port, 
      fifo_0_8_port, fifo_0_7_port, fifo_0_6_port, fifo_0_5_port, fifo_0_4_port
      , fifo_0_3_port, fifo_0_2_port, fifo_0_1_port, fifo_0_0_port, N7, N9, n1,
      n3, n5, n7_port, n9_port, n11, n13, n15, n17, n19, n21, n23, n25, n27, 
      n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57
      , n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, 
      n87, n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, n111, 
      n113, n115, n117, n119, n121, n123, n125, n127, n129, n131, n133, n135, 
      n137, n139, n141, n143, n145, n147, n149, n151, n153, n155, n157, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238 : std_logic;

begin
   valid_data <= valid_data_port;
   
   U4 : XOR2xp5_ASAP7_75t_R port map( A => N7, B => n43, Y => n238);
   U143 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_9_port, B1 => 
                           n43, B2 => fifo_0_9_port, Y => data_out(9));
   U144 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_8_port, B1 => 
                           n43, B2 => fifo_0_8_port, Y => data_out(8));
   U145 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_7_port, B1 => 
                           n43, B2 => fifo_0_7_port, Y => data_out(7));
   U146 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_6_port, B1 => 
                           n43, B2 => fifo_0_6_port, Y => data_out(6));
   U147 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_63_port, B1 => 
                           n43, B2 => fifo_0_63_port, Y => data_out(63));
   U148 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_62_port, B1 => 
                           n43, B2 => fifo_0_62_port, Y => data_out(62));
   U149 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_61_port, B1 => 
                           n43, B2 => fifo_0_61_port, Y => data_out(61));
   U150 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_60_port, B1 => 
                           n43, B2 => fifo_0_60_port, Y => data_out(60));
   U151 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_5_port, B1 => 
                           n43, B2 => fifo_0_5_port, Y => data_out(5));
   U152 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_59_port, B1 => 
                           n43, B2 => fifo_0_59_port, Y => data_out(59));
   U153 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_58_port, B1 => 
                           n43, B2 => fifo_0_58_port, Y => data_out(58));
   U154 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_57_port, B1 => 
                           n43, B2 => fifo_0_57_port, Y => data_out(57));
   U155 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_56_port, B1 => 
                           n43, B2 => fifo_0_56_port, Y => data_out(56));
   U156 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_55_port, B1 => 
                           n43, B2 => fifo_0_55_port, Y => data_out(55));
   U157 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_54_port, B1 => 
                           n43, B2 => fifo_0_54_port, Y => data_out(54));
   U158 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_53_port, B1 => 
                           n43, B2 => fifo_0_53_port, Y => data_out(53));
   U159 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_52_port, B1 => 
                           n43, B2 => fifo_0_52_port, Y => data_out(52));
   U160 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_51_port, B1 => 
                           n43, B2 => fifo_0_51_port, Y => data_out(51));
   U161 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_50_port, B1 => 
                           n43, B2 => fifo_0_50_port, Y => data_out(50));
   U162 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_4_port, B1 => 
                           n43, B2 => fifo_0_4_port, Y => data_out(4));
   U163 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_49_port, B1 => 
                           n43, B2 => fifo_0_49_port, Y => data_out(49));
   U164 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_48_port, B1 => 
                           n43, B2 => fifo_0_48_port, Y => data_out(48));
   U165 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_47_port, B1 => 
                           n43, B2 => fifo_0_47_port, Y => data_out(47));
   U166 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_46_port, B1 => 
                           n43, B2 => fifo_0_46_port, Y => data_out(46));
   U167 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_45_port, B1 => 
                           n43, B2 => fifo_0_45_port, Y => data_out(45));
   U168 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_44_port, B1 => 
                           n43, B2 => fifo_0_44_port, Y => data_out(44));
   U169 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_43_port, B1 => 
                           n43, B2 => fifo_0_43_port, Y => data_out(43));
   U170 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_42_port, B1 => 
                           n43, B2 => fifo_0_42_port, Y => data_out(42));
   U171 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_41_port, B1 => 
                           n43, B2 => fifo_0_41_port, Y => data_out(41));
   U172 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_40_port, B1 => 
                           n43, B2 => fifo_0_40_port, Y => data_out(40));
   U173 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_3_port, B1 => 
                           n43, B2 => fifo_0_3_port, Y => data_out(3));
   U174 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_39_port, B1 => 
                           n43, B2 => fifo_0_39_port, Y => data_out(39));
   U175 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_38_port, B1 => 
                           n43, B2 => fifo_0_38_port, Y => data_out(38));
   U176 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_37_port, B1 => 
                           n43, B2 => fifo_0_37_port, Y => data_out(37));
   U177 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_36_port, B1 => 
                           n43, B2 => fifo_0_36_port, Y => data_out(36));
   U178 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_35_port, B1 => 
                           n43, B2 => fifo_0_35_port, Y => data_out(35));
   U179 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_34_port, B1 => 
                           n43, B2 => fifo_0_34_port, Y => data_out(34));
   U180 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_33_port, B1 => 
                           n43, B2 => fifo_0_33_port, Y => data_out(33));
   U181 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_32_port, B1 => 
                           n43, B2 => fifo_0_32_port, Y => data_out(32));
   U182 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_31_port, B1 => 
                           n43, B2 => fifo_0_31_port, Y => data_out(31));
   U183 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_30_port, B1 => 
                           n43, B2 => fifo_0_30_port, Y => data_out(30));
   U184 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_2_port, B1 => 
                           n43, B2 => fifo_0_2_port, Y => data_out(2));
   U185 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_29_port, B1 => 
                           n43, B2 => fifo_0_29_port, Y => data_out(29));
   U186 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_28_port, B1 => 
                           n43, B2 => fifo_0_28_port, Y => data_out(28));
   U187 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_27_port, B1 => 
                           n43, B2 => fifo_0_27_port, Y => data_out(27));
   U188 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_26_port, B1 => 
                           n43, B2 => fifo_0_26_port, Y => data_out(26));
   U189 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_25_port, B1 => 
                           n43, B2 => fifo_0_25_port, Y => data_out(25));
   U190 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_24_port, B1 => 
                           n43, B2 => fifo_0_24_port, Y => data_out(24));
   U191 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_23_port, B1 => 
                           n43, B2 => fifo_0_23_port, Y => data_out(23));
   U192 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_22_port, B1 => 
                           n43, B2 => fifo_0_22_port, Y => data_out(22));
   U193 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_21_port, B1 => 
                           n43, B2 => fifo_0_21_port, Y => data_out(21));
   U194 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_20_port, B1 => 
                           n43, B2 => fifo_0_20_port, Y => data_out(20));
   U195 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_1_port, B1 => 
                           n43, B2 => fifo_0_1_port, Y => data_out(1));
   U196 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_19_port, B1 => 
                           n43, B2 => fifo_0_19_port, Y => data_out(19));
   U197 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_18_port, B1 => 
                           n43, B2 => fifo_0_18_port, Y => data_out(18));
   U198 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_17_port, B1 => 
                           n43, B2 => fifo_0_17_port, Y => data_out(17));
   U199 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_16_port, B1 => 
                           n43, B2 => fifo_0_16_port, Y => data_out(16));
   U200 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_15_port, B1 => 
                           n43, B2 => fifo_0_15_port, Y => data_out(15));
   U201 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_14_port, B1 => 
                           n43, B2 => fifo_0_14_port, Y => data_out(14));
   U202 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_13_port, B1 => 
                           n43, B2 => fifo_0_13_port, Y => data_out(13));
   U203 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_12_port, B1 => 
                           n43, B2 => fifo_0_12_port, Y => data_out(12));
   U204 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_11_port, B1 => 
                           n43, B2 => fifo_0_11_port, Y => data_out(11));
   U205 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_10_port, B1 => 
                           n43, B2 => fifo_0_10_port, Y => data_out(10));
   U206 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_0_port, B1 => 
                           n43, B2 => fifo_0_0_port, Y => data_out(0));
   U3 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n45, A2 => n238, B => 
                           valid_data_port, C => write_en, Y => n235);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_0_port, A2 => n17, B1 => 
                           data_in(0), B2 => n29, Y => n234);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_1_port, A2 => n17, B1 => 
                           data_in(1), B2 => n29, Y => n233);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_2_port, A2 => n17, B1 => 
                           data_in(2), B2 => n29, Y => n232);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_3_port, A2 => n17, B1 => 
                           data_in(3), B2 => n29, Y => n231);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_4_port, A2 => n17, B1 => 
                           data_in(4), B2 => n27, Y => n230);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_5_port, A2 => n17, B1 => 
                           data_in(5), B2 => n27, Y => n229);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_6_port, A2 => n17, B1 => 
                           data_in(6), B2 => n27, Y => n228);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_7_port, A2 => n17, B1 => 
                           data_in(7), B2 => n27, Y => n227);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_8_port, A2 => n17, B1 => 
                           data_in(8), B2 => n27, Y => n226);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_9_port, A2 => n17, B1 => 
                           data_in(9), B2 => n27, Y => n225);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_10_port, A2 => n17, B1 => 
                           data_in(10), B2 => n27, Y => n224);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_11_port, A2 => n17, B1 => 
                           data_in(11), B2 => n27, Y => n223);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_12_port, A2 => n17, B1 => 
                           data_in(12), B2 => n27, Y => n222);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_13_port, A2 => n17, B1 => 
                           data_in(13), B2 => n27, Y => n221);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_14_port, A2 => n17, B1 => 
                           data_in(14), B2 => n27, Y => n220);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_15_port, A2 => n17, B1 => 
                           data_in(15), B2 => n27, Y => n219);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_16_port, A2 => n17, B1 => 
                           data_in(16), B2 => n25, Y => n218);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_17_port, A2 => n17, B1 => 
                           data_in(17), B2 => n25, Y => n217);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_18_port, A2 => n17, B1 => 
                           data_in(18), B2 => n25, Y => n216);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_19_port, A2 => n17, B1 => 
                           data_in(19), B2 => n25, Y => n215);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_20_port, A2 => n17, B1 => 
                           data_in(20), B2 => n25, Y => n214);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_21_port, A2 => n17, B1 => 
                           data_in(21), B2 => n25, Y => n213);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_22_port, A2 => n17, B1 => 
                           data_in(22), B2 => n25, Y => n212);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_23_port, A2 => n17, B1 => 
                           data_in(23), B2 => n25, Y => n211);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_24_port, A2 => n17, B1 => 
                           data_in(24), B2 => n25, Y => n210);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_25_port, A2 => n17, B1 => 
                           data_in(25), B2 => n25, Y => n209);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_26_port, A2 => n17, B1 => 
                           data_in(26), B2 => n25, Y => n208);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_27_port, A2 => n17, B1 => 
                           data_in(27), B2 => n25, Y => n207);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_28_port, A2 => n17, B1 => 
                           data_in(28), B2 => n23, Y => n206);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_29_port, A2 => n17, B1 => 
                           data_in(29), B2 => n23, Y => n205);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_30_port, A2 => n17, B1 => 
                           data_in(30), B2 => n23, Y => n204);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_31_port, A2 => n17, B1 => 
                           data_in(31), B2 => n23, Y => n203);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_32_port, A2 => n17, B1 => 
                           data_in(32), B2 => n23, Y => n202);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_33_port, A2 => n17, B1 => 
                           data_in(33), B2 => n23, Y => n201);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_34_port, A2 => n17, B1 => 
                           data_in(34), B2 => n23, Y => n200);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_35_port, A2 => n17, B1 => 
                           data_in(35), B2 => n23, Y => n199);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_36_port, A2 => n17, B1 => 
                           data_in(36), B2 => n23, Y => n198);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_37_port, A2 => n17, B1 => 
                           data_in(37), B2 => n23, Y => n197);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_38_port, A2 => n17, B1 => 
                           data_in(38), B2 => n23, Y => n196);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_39_port, A2 => n17, B1 => 
                           data_in(39), B2 => n23, Y => n195);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_40_port, A2 => n17, B1 => 
                           data_in(40), B2 => n21, Y => n194);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_41_port, A2 => n17, B1 => 
                           data_in(41), B2 => n21, Y => n193);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_42_port, A2 => n17, B1 => 
                           data_in(42), B2 => n21, Y => n192);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_43_port, A2 => n17, B1 => 
                           data_in(43), B2 => n21, Y => n191);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_44_port, A2 => n17, B1 => 
                           data_in(44), B2 => n21, Y => n190);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_45_port, A2 => n17, B1 => 
                           data_in(45), B2 => n21, Y => n189);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_46_port, A2 => n17, B1 => 
                           data_in(46), B2 => n21, Y => n188);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_47_port, A2 => n17, B1 => 
                           data_in(47), B2 => n21, Y => n187);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_48_port, A2 => n17, B1 => 
                           data_in(48), B2 => n21, Y => n186);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_49_port, A2 => n17, B1 => 
                           data_in(49), B2 => n21, Y => n185);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_50_port, A2 => n17, B1 => 
                           data_in(50), B2 => n21, Y => n184);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_51_port, A2 => n17, B1 => 
                           data_in(51), B2 => n21, Y => n183);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_52_port, A2 => n17, B1 => 
                           data_in(52), B2 => n19, Y => n182);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_53_port, A2 => n17, B1 => 
                           data_in(53), B2 => n19, Y => n181);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_54_port, A2 => n17, B1 => 
                           data_in(54), B2 => n19, Y => n180);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_55_port, A2 => n17, B1 => 
                           data_in(55), B2 => n19, Y => n179);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_56_port, A2 => n17, B1 => 
                           data_in(56), B2 => n19, Y => n178);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_57_port, A2 => n17, B1 => 
                           data_in(57), B2 => n19, Y => n177);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_58_port, A2 => n17, B1 => 
                           data_in(58), B2 => n19, Y => n176);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_59_port, A2 => n17, B1 => 
                           data_in(59), B2 => n19, Y => n175);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_60_port, A2 => n17, B1 => 
                           data_in(60), B2 => n19, Y => n174);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_61_port, A2 => n17, B1 => 
                           data_in(61), B2 => n19, Y => n173);
   U67 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_62_port, A2 => n17, B1 => 
                           data_in(62), B2 => n19, Y => n172);
   U68 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_63_port, A2 => n17, B1 => 
                           data_in(63), B2 => n19, Y => n171);
   U70 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N9, Y => n237);
   U71 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_0_port, A2 => n3, B1 => 
                           data_in(0), B2 => n15, Y => n170);
   U72 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_1_port, A2 => n3, B1 => 
                           data_in(1), B2 => n15, Y => n169);
   U73 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_2_port, A2 => n3, B1 => 
                           data_in(2), B2 => n15, Y => n168);
   U74 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_3_port, A2 => n3, B1 => 
                           data_in(3), B2 => n15, Y => n167);
   U75 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_4_port, A2 => n3, B1 => 
                           data_in(4), B2 => n13, Y => n166);
   U76 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_5_port, A2 => n3, B1 => 
                           data_in(5), B2 => n13, Y => n165);
   U77 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_6_port, A2 => n3, B1 => 
                           data_in(6), B2 => n13, Y => n164);
   U78 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_7_port, A2 => n3, B1 => 
                           data_in(7), B2 => n13, Y => n163);
   U79 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_8_port, A2 => n3, B1 => 
                           data_in(8), B2 => n13, Y => n162);
   U80 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_9_port, A2 => n3, B1 => 
                           data_in(9), B2 => n13, Y => n161);
   U81 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_10_port, A2 => n3, B1 => 
                           data_in(10), B2 => n13, Y => n160);
   U82 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_11_port, A2 => n3, B1 => 
                           data_in(11), B2 => n13, Y => n159);
   U83 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_12_port, A2 => n3, B1 => 
                           data_in(12), B2 => n13, Y => n157);
   U84 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_13_port, A2 => n3, B1 => 
                           data_in(13), B2 => n13, Y => n155);
   U85 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_14_port, A2 => n3, B1 => 
                           data_in(14), B2 => n13, Y => n153);
   U86 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_15_port, A2 => n3, B1 => 
                           data_in(15), B2 => n13, Y => n151);
   U87 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_16_port, A2 => n3, B1 => 
                           data_in(16), B2 => n11, Y => n149);
   U88 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_17_port, A2 => n3, B1 => 
                           data_in(17), B2 => n11, Y => n147);
   U89 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_18_port, A2 => n3, B1 => 
                           data_in(18), B2 => n11, Y => n145);
   U90 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_19_port, A2 => n3, B1 => 
                           data_in(19), B2 => n11, Y => n143);
   U91 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_20_port, A2 => n3, B1 => 
                           data_in(20), B2 => n11, Y => n141);
   U92 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_21_port, A2 => n3, B1 => 
                           data_in(21), B2 => n11, Y => n139);
   U93 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_22_port, A2 => n3, B1 => 
                           data_in(22), B2 => n11, Y => n137);
   U94 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_23_port, A2 => n3, B1 => 
                           data_in(23), B2 => n11, Y => n135);
   U95 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_24_port, A2 => n3, B1 => 
                           data_in(24), B2 => n11, Y => n133);
   U96 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_25_port, A2 => n3, B1 => 
                           data_in(25), B2 => n11, Y => n131);
   U97 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_26_port, A2 => n3, B1 => 
                           data_in(26), B2 => n11, Y => n129);
   U98 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_27_port, A2 => n3, B1 => 
                           data_in(27), B2 => n11, Y => n127);
   U99 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_28_port, A2 => n3, B1 => 
                           data_in(28), B2 => n9_port, Y => n125);
   U100 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_29_port, A2 => n3, B1 => 
                           data_in(29), B2 => n9_port, Y => n123);
   U101 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_30_port, A2 => n3, B1 => 
                           data_in(30), B2 => n9_port, Y => n121);
   U102 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_31_port, A2 => n3, B1 => 
                           data_in(31), B2 => n9_port, Y => n119);
   U103 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_32_port, A2 => n3, B1 => 
                           data_in(32), B2 => n9_port, Y => n117);
   U104 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_33_port, A2 => n3, B1 => 
                           data_in(33), B2 => n9_port, Y => n115);
   U105 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_34_port, A2 => n3, B1 => 
                           data_in(34), B2 => n9_port, Y => n113);
   U106 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_35_port, A2 => n3, B1 => 
                           data_in(35), B2 => n9_port, Y => n111);
   U107 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_36_port, A2 => n3, B1 => 
                           data_in(36), B2 => n9_port, Y => n109);
   U108 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_37_port, A2 => n3, B1 => 
                           data_in(37), B2 => n9_port, Y => n107);
   U109 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_38_port, A2 => n3, B1 => 
                           data_in(38), B2 => n9_port, Y => n105);
   U110 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_39_port, A2 => n3, B1 => 
                           data_in(39), B2 => n9_port, Y => n103);
   U111 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_40_port, A2 => n3, B1 => 
                           data_in(40), B2 => n7_port, Y => n101);
   U112 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_41_port, A2 => n3, B1 => 
                           data_in(41), B2 => n7_port, Y => n99);
   U113 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_42_port, A2 => n3, B1 => 
                           data_in(42), B2 => n7_port, Y => n97);
   U114 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_43_port, A2 => n3, B1 => 
                           data_in(43), B2 => n7_port, Y => n95);
   U115 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_44_port, A2 => n3, B1 => 
                           data_in(44), B2 => n7_port, Y => n93);
   U116 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_45_port, A2 => n3, B1 => 
                           data_in(45), B2 => n7_port, Y => n91);
   U117 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_46_port, A2 => n3, B1 => 
                           data_in(46), B2 => n7_port, Y => n89);
   U118 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_47_port, A2 => n3, B1 => 
                           data_in(47), B2 => n7_port, Y => n87);
   U119 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_48_port, A2 => n3, B1 => 
                           data_in(48), B2 => n7_port, Y => n85);
   U120 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_49_port, A2 => n3, B1 => 
                           data_in(49), B2 => n7_port, Y => n83);
   U121 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_50_port, A2 => n3, B1 => 
                           data_in(50), B2 => n7_port, Y => n81);
   U122 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_51_port, A2 => n3, B1 => 
                           data_in(51), B2 => n7_port, Y => n79);
   U123 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_52_port, A2 => n3, B1 => 
                           data_in(52), B2 => n5, Y => n77);
   U124 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_53_port, A2 => n3, B1 => 
                           data_in(53), B2 => n5, Y => n75);
   U125 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_54_port, A2 => n3, B1 => 
                           data_in(54), B2 => n5, Y => n73);
   U126 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_55_port, A2 => n3, B1 => 
                           data_in(55), B2 => n5, Y => n71);
   U127 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_56_port, A2 => n3, B1 => 
                           data_in(56), B2 => n5, Y => n69);
   U128 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_57_port, A2 => n3, B1 => 
                           data_in(57), B2 => n5, Y => n67);
   U129 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_58_port, A2 => n3, B1 => 
                           data_in(58), B2 => n5, Y => n65);
   U130 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_59_port, A2 => n3, B1 => 
                           data_in(59), B2 => n5, Y => n63);
   U131 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_60_port, A2 => n3, B1 => 
                           data_in(60), B2 => n5, Y => n61);
   U132 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_61_port, A2 => n3, B1 => 
                           data_in(61), B2 => n5, Y => n59);
   U133 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_62_port, A2 => n3, B1 => 
                           data_in(62), B2 => n5, Y => n57);
   U134 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_63_port, A2 => n3, B1 => 
                           data_in(63), B2 => n5, Y => n55);
   U136 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N7, Y => n236);
   U137 : OAI22xp5_ASAP7_75t_R port map( A1 => n31, A2 => read_en, B1 => n43, 
                           B2 => n45, Y => n53);
   U139 : OAI22xp5_ASAP7_75t_R port map( A1 => N9, A2 => n49, B1 => write_en, 
                           B2 => N7, Y => n51);
   write_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK 
                           => clk, RESET => n47, SET => n1, QN => N7);
   fifo_reg_1_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n55, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_63_port);
   fifo_reg_1_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n57, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_62_port);
   fifo_reg_1_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n59, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_61_port);
   fifo_reg_1_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n61, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_60_port);
   fifo_reg_0_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n171, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_63_port);
   fifo_reg_0_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n172, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_62_port);
   fifo_reg_0_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n173, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_61_port);
   fifo_reg_0_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n174, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_60_port);
   fifo_reg_1_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n167, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_3_port);
   fifo_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n168, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_2_port);
   fifo_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n169, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_1_port);
   fifo_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n170, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_0_port);
   fifo_reg_1_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n63, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_59_port);
   fifo_reg_1_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n65, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_58_port);
   fifo_reg_1_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n67, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_57_port);
   fifo_reg_1_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n69, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_56_port);
   fifo_reg_1_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n71, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_55_port);
   fifo_reg_1_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n73, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_54_port);
   fifo_reg_1_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n75, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_53_port);
   fifo_reg_1_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n77, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_52_port);
   fifo_reg_1_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_51_port);
   fifo_reg_1_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_50_port);
   fifo_reg_1_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_49_port);
   fifo_reg_1_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_48_port);
   fifo_reg_1_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_47_port);
   fifo_reg_1_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_46_port);
   fifo_reg_1_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_45_port);
   fifo_reg_1_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_44_port);
   fifo_reg_1_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_43_port);
   fifo_reg_1_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_42_port);
   fifo_reg_1_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_41_port);
   fifo_reg_1_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_40_port);
   fifo_reg_1_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_39_port);
   fifo_reg_1_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_38_port);
   fifo_reg_1_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_37_port);
   fifo_reg_1_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_36_port);
   fifo_reg_1_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_35_port);
   fifo_reg_1_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_34_port);
   fifo_reg_1_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n115, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_33_port);
   fifo_reg_1_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n117, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_32_port);
   fifo_reg_1_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n119, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_31_port);
   fifo_reg_1_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n121, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_30_port);
   fifo_reg_1_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n123, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_29_port);
   fifo_reg_1_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n125, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_28_port);
   fifo_reg_1_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n127, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_27_port);
   fifo_reg_1_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n129, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_26_port);
   fifo_reg_1_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n131, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_25_port);
   fifo_reg_1_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n133, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_24_port);
   fifo_reg_1_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n135, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_23_port);
   fifo_reg_1_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n137, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_22_port);
   fifo_reg_1_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n139, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_21_port);
   fifo_reg_1_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n141, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_20_port);
   fifo_reg_1_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n143, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_19_port);
   fifo_reg_1_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n145, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_18_port);
   fifo_reg_1_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n147, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_17_port);
   fifo_reg_1_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n149, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_16_port);
   fifo_reg_1_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n151, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_15_port);
   fifo_reg_1_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n153, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_14_port);
   fifo_reg_1_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n155, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_13_port);
   fifo_reg_1_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n157, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_12_port);
   fifo_reg_1_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n159, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_11_port);
   fifo_reg_1_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n160, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_10_port);
   fifo_reg_1_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n161, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_9_port);
   fifo_reg_1_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n162, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_8_port);
   fifo_reg_1_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n163, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_7_port);
   fifo_reg_1_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n164, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_6_port);
   fifo_reg_1_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n165, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_5_port);
   fifo_reg_1_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n166, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_4_port);
   fifo_reg_0_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n231, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_3_port);
   fifo_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n232, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_2_port);
   fifo_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n233, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_1_port);
   fifo_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n234, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_0_port);
   fifo_reg_0_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n175, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_59_port);
   fifo_reg_0_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n176, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_58_port);
   fifo_reg_0_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n177, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_57_port);
   fifo_reg_0_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n178, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_56_port);
   fifo_reg_0_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n179, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_55_port);
   fifo_reg_0_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n180, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_54_port);
   fifo_reg_0_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n181, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_53_port);
   fifo_reg_0_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n182, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_52_port);
   fifo_reg_0_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n183, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_51_port);
   fifo_reg_0_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n184, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_50_port);
   fifo_reg_0_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n185, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_49_port);
   fifo_reg_0_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n186, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_48_port);
   fifo_reg_0_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n187, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_47_port);
   fifo_reg_0_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n188, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_46_port);
   fifo_reg_0_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n189, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_45_port);
   fifo_reg_0_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n190, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_44_port);
   fifo_reg_0_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n191, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_43_port);
   fifo_reg_0_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n192, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_42_port);
   fifo_reg_0_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n193, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_41_port);
   fifo_reg_0_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n194, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_40_port);
   fifo_reg_0_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n195, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_39_port);
   fifo_reg_0_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n196, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_38_port);
   fifo_reg_0_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n197, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_37_port);
   fifo_reg_0_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n198, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_36_port);
   fifo_reg_0_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n199, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_35_port);
   fifo_reg_0_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n200, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_34_port);
   fifo_reg_0_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n201, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_33_port);
   fifo_reg_0_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n202, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_32_port);
   fifo_reg_0_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n203, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_31_port);
   fifo_reg_0_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n204, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_30_port);
   fifo_reg_0_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n205, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_29_port);
   fifo_reg_0_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n206, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_28_port);
   fifo_reg_0_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n207, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_27_port);
   fifo_reg_0_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n208, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_26_port);
   fifo_reg_0_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n209, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_25_port);
   fifo_reg_0_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n210, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_24_port);
   fifo_reg_0_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n211, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_23_port);
   fifo_reg_0_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n212, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_22_port);
   fifo_reg_0_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n213, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_21_port);
   fifo_reg_0_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n214, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_20_port);
   fifo_reg_0_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n215, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_19_port);
   fifo_reg_0_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n216, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_18_port);
   fifo_reg_0_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n217, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_17_port);
   fifo_reg_0_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n218, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_16_port);
   fifo_reg_0_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n219, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_15_port);
   fifo_reg_0_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n220, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_14_port);
   fifo_reg_0_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n221, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_13_port);
   fifo_reg_0_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n222, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_12_port);
   fifo_reg_0_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n223, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_11_port);
   fifo_reg_0_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n224, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_10_port);
   fifo_reg_0_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n225, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_9_port);
   fifo_reg_0_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n226, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_8_port);
   fifo_reg_0_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n227, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_7_port);
   fifo_reg_0_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n228, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_6_port);
   fifo_reg_0_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n229, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_5_port);
   fifo_reg_0_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n230, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_4_port);
   valid_data_reg : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n235, CLK => clk, 
                           RESET => n47, SET => n1, QN => valid_data_port);
   read_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK 
                           => clk, RESET => n47, SET => n1, QN => 
                           read_pointer_0_port);
   U69 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U135 : INVx3_ASAP7_75t_R port map( A => rst, Y => n47);
   U138 : INVx1_ASAP7_75t_R port map( A => read_en, Y => n45);
   U140 : INVx1_ASAP7_75t_R port map( A => n29, Y => n17);
   U141 : INVx1_ASAP7_75t_R port map( A => n15, Y => n3);
   U142 : INVx1_ASAP7_75t_R port map( A => n31, Y => n43);
   U207 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n29);
   U208 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n15);
   U209 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n27);
   U210 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n25);
   U211 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n23);
   U212 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n21);
   U213 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n19);
   U214 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n13);
   U215 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n11);
   U216 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n9_port);
   U217 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n7_port);
   U218 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n5);
   U219 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n31);
   U220 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n33);
   U221 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n41);
   U222 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n39);
   U223 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n37);
   U224 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n35);
   U225 : INVx1_ASAP7_75t_R port map( A => N7, Y => N9);
   U226 : INVx1_ASAP7_75t_R port map( A => write_en, Y => n49);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity fifo_buff_depth2_4 is

   port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, clk, 
         rst : in std_logic;  data_out : out std_logic_vector (63 downto 0);  
         valid_data : out std_logic);

end fifo_buff_depth2_4;

architecture SYN_rtl of fifo_buff_depth2_4 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx3_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal valid_data_port, read_pointer_0_port, fifo_1_63_port, fifo_1_62_port,
      fifo_1_61_port, fifo_1_60_port, fifo_1_59_port, fifo_1_58_port, 
      fifo_1_57_port, fifo_1_56_port, fifo_1_55_port, fifo_1_54_port, 
      fifo_1_53_port, fifo_1_52_port, fifo_1_51_port, fifo_1_50_port, 
      fifo_1_49_port, fifo_1_48_port, fifo_1_47_port, fifo_1_46_port, 
      fifo_1_45_port, fifo_1_44_port, fifo_1_43_port, fifo_1_42_port, 
      fifo_1_41_port, fifo_1_40_port, fifo_1_39_port, fifo_1_38_port, 
      fifo_1_37_port, fifo_1_36_port, fifo_1_35_port, fifo_1_34_port, 
      fifo_1_33_port, fifo_1_32_port, fifo_1_31_port, fifo_1_30_port, 
      fifo_1_29_port, fifo_1_28_port, fifo_1_27_port, fifo_1_26_port, 
      fifo_1_25_port, fifo_1_24_port, fifo_1_23_port, fifo_1_22_port, 
      fifo_1_21_port, fifo_1_20_port, fifo_1_19_port, fifo_1_18_port, 
      fifo_1_17_port, fifo_1_16_port, fifo_1_15_port, fifo_1_14_port, 
      fifo_1_13_port, fifo_1_12_port, fifo_1_11_port, fifo_1_10_port, 
      fifo_1_9_port, fifo_1_8_port, fifo_1_7_port, fifo_1_6_port, fifo_1_5_port
      , fifo_1_4_port, fifo_1_3_port, fifo_1_2_port, fifo_1_1_port, 
      fifo_1_0_port, fifo_0_63_port, fifo_0_62_port, fifo_0_61_port, 
      fifo_0_60_port, fifo_0_59_port, fifo_0_58_port, fifo_0_57_port, 
      fifo_0_56_port, fifo_0_55_port, fifo_0_54_port, fifo_0_53_port, 
      fifo_0_52_port, fifo_0_51_port, fifo_0_50_port, fifo_0_49_port, 
      fifo_0_48_port, fifo_0_47_port, fifo_0_46_port, fifo_0_45_port, 
      fifo_0_44_port, fifo_0_43_port, fifo_0_42_port, fifo_0_41_port, 
      fifo_0_40_port, fifo_0_39_port, fifo_0_38_port, fifo_0_37_port, 
      fifo_0_36_port, fifo_0_35_port, fifo_0_34_port, fifo_0_33_port, 
      fifo_0_32_port, fifo_0_31_port, fifo_0_30_port, fifo_0_29_port, 
      fifo_0_28_port, fifo_0_27_port, fifo_0_26_port, fifo_0_25_port, 
      fifo_0_24_port, fifo_0_23_port, fifo_0_22_port, fifo_0_21_port, 
      fifo_0_20_port, fifo_0_19_port, fifo_0_18_port, fifo_0_17_port, 
      fifo_0_16_port, fifo_0_15_port, fifo_0_14_port, fifo_0_13_port, 
      fifo_0_12_port, fifo_0_11_port, fifo_0_10_port, fifo_0_9_port, 
      fifo_0_8_port, fifo_0_7_port, fifo_0_6_port, fifo_0_5_port, fifo_0_4_port
      , fifo_0_3_port, fifo_0_2_port, fifo_0_1_port, fifo_0_0_port, N7, N9, n1,
      n3, n5, n7_port, n9_port, n11, n13, n15, n17, n19, n21, n23, n25, n27, 
      n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57
      , n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, 
      n87, n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, n111, 
      n113, n115, n117, n119, n121, n123, n125, n127, n129, n131, n133, n135, 
      n137, n139, n141, n143, n145, n147, n149, n151, n153, n155, n157, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238 : std_logic;

begin
   valid_data <= valid_data_port;
   
   U4 : XOR2xp5_ASAP7_75t_R port map( A => N7, B => n43, Y => n238);
   U143 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_9_port, B1 => 
                           n43, B2 => fifo_0_9_port, Y => data_out(9));
   U144 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_8_port, B1 => 
                           n43, B2 => fifo_0_8_port, Y => data_out(8));
   U145 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_7_port, B1 => 
                           n43, B2 => fifo_0_7_port, Y => data_out(7));
   U146 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_6_port, B1 => 
                           n43, B2 => fifo_0_6_port, Y => data_out(6));
   U147 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_63_port, B1 => 
                           n43, B2 => fifo_0_63_port, Y => data_out(63));
   U148 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_62_port, B1 => 
                           n43, B2 => fifo_0_62_port, Y => data_out(62));
   U149 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_61_port, B1 => 
                           n43, B2 => fifo_0_61_port, Y => data_out(61));
   U150 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_60_port, B1 => 
                           n43, B2 => fifo_0_60_port, Y => data_out(60));
   U151 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_5_port, B1 => 
                           n43, B2 => fifo_0_5_port, Y => data_out(5));
   U152 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_59_port, B1 => 
                           n43, B2 => fifo_0_59_port, Y => data_out(59));
   U153 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_58_port, B1 => 
                           n43, B2 => fifo_0_58_port, Y => data_out(58));
   U154 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_57_port, B1 => 
                           n43, B2 => fifo_0_57_port, Y => data_out(57));
   U155 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_56_port, B1 => 
                           n43, B2 => fifo_0_56_port, Y => data_out(56));
   U156 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_55_port, B1 => 
                           n43, B2 => fifo_0_55_port, Y => data_out(55));
   U157 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_54_port, B1 => 
                           n43, B2 => fifo_0_54_port, Y => data_out(54));
   U158 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_53_port, B1 => 
                           n43, B2 => fifo_0_53_port, Y => data_out(53));
   U159 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_52_port, B1 => 
                           n43, B2 => fifo_0_52_port, Y => data_out(52));
   U160 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_51_port, B1 => 
                           n43, B2 => fifo_0_51_port, Y => data_out(51));
   U161 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_50_port, B1 => 
                           n43, B2 => fifo_0_50_port, Y => data_out(50));
   U162 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_4_port, B1 => 
                           n43, B2 => fifo_0_4_port, Y => data_out(4));
   U163 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_49_port, B1 => 
                           n43, B2 => fifo_0_49_port, Y => data_out(49));
   U164 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_48_port, B1 => 
                           n43, B2 => fifo_0_48_port, Y => data_out(48));
   U165 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_47_port, B1 => 
                           n43, B2 => fifo_0_47_port, Y => data_out(47));
   U166 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_46_port, B1 => 
                           n43, B2 => fifo_0_46_port, Y => data_out(46));
   U167 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_45_port, B1 => 
                           n43, B2 => fifo_0_45_port, Y => data_out(45));
   U168 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_44_port, B1 => 
                           n43, B2 => fifo_0_44_port, Y => data_out(44));
   U169 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_43_port, B1 => 
                           n43, B2 => fifo_0_43_port, Y => data_out(43));
   U170 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_42_port, B1 => 
                           n43, B2 => fifo_0_42_port, Y => data_out(42));
   U171 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_41_port, B1 => 
                           n43, B2 => fifo_0_41_port, Y => data_out(41));
   U172 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_40_port, B1 => 
                           n43, B2 => fifo_0_40_port, Y => data_out(40));
   U173 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_3_port, B1 => 
                           n43, B2 => fifo_0_3_port, Y => data_out(3));
   U174 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_39_port, B1 => 
                           n43, B2 => fifo_0_39_port, Y => data_out(39));
   U175 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_38_port, B1 => 
                           n43, B2 => fifo_0_38_port, Y => data_out(38));
   U176 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_37_port, B1 => 
                           n43, B2 => fifo_0_37_port, Y => data_out(37));
   U177 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_36_port, B1 => 
                           n43, B2 => fifo_0_36_port, Y => data_out(36));
   U178 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_35_port, B1 => 
                           n43, B2 => fifo_0_35_port, Y => data_out(35));
   U179 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_34_port, B1 => 
                           n43, B2 => fifo_0_34_port, Y => data_out(34));
   U180 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_33_port, B1 => 
                           n43, B2 => fifo_0_33_port, Y => data_out(33));
   U181 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_32_port, B1 => 
                           n43, B2 => fifo_0_32_port, Y => data_out(32));
   U182 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_31_port, B1 => 
                           n43, B2 => fifo_0_31_port, Y => data_out(31));
   U183 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_30_port, B1 => 
                           n43, B2 => fifo_0_30_port, Y => data_out(30));
   U184 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_2_port, B1 => 
                           n43, B2 => fifo_0_2_port, Y => data_out(2));
   U185 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_29_port, B1 => 
                           n43, B2 => fifo_0_29_port, Y => data_out(29));
   U186 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_28_port, B1 => 
                           n43, B2 => fifo_0_28_port, Y => data_out(28));
   U187 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_27_port, B1 => 
                           n43, B2 => fifo_0_27_port, Y => data_out(27));
   U188 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_26_port, B1 => 
                           n43, B2 => fifo_0_26_port, Y => data_out(26));
   U189 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_25_port, B1 => 
                           n43, B2 => fifo_0_25_port, Y => data_out(25));
   U190 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_24_port, B1 => 
                           n43, B2 => fifo_0_24_port, Y => data_out(24));
   U191 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_23_port, B1 => 
                           n43, B2 => fifo_0_23_port, Y => data_out(23));
   U192 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_22_port, B1 => 
                           n43, B2 => fifo_0_22_port, Y => data_out(22));
   U193 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_21_port, B1 => 
                           n43, B2 => fifo_0_21_port, Y => data_out(21));
   U194 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_20_port, B1 => 
                           n43, B2 => fifo_0_20_port, Y => data_out(20));
   U195 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_1_port, B1 => 
                           n43, B2 => fifo_0_1_port, Y => data_out(1));
   U196 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_19_port, B1 => 
                           n43, B2 => fifo_0_19_port, Y => data_out(19));
   U197 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_18_port, B1 => 
                           n43, B2 => fifo_0_18_port, Y => data_out(18));
   U198 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_17_port, B1 => 
                           n43, B2 => fifo_0_17_port, Y => data_out(17));
   U199 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_16_port, B1 => 
                           n43, B2 => fifo_0_16_port, Y => data_out(16));
   U200 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_15_port, B1 => 
                           n43, B2 => fifo_0_15_port, Y => data_out(15));
   U201 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_14_port, B1 => 
                           n43, B2 => fifo_0_14_port, Y => data_out(14));
   U202 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_13_port, B1 => 
                           n43, B2 => fifo_0_13_port, Y => data_out(13));
   U203 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_12_port, B1 => 
                           n43, B2 => fifo_0_12_port, Y => data_out(12));
   U204 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_11_port, B1 => 
                           n43, B2 => fifo_0_11_port, Y => data_out(11));
   U205 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_10_port, B1 => 
                           n43, B2 => fifo_0_10_port, Y => data_out(10));
   U206 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_0_port, B1 => 
                           n43, B2 => fifo_0_0_port, Y => data_out(0));
   U3 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n47, A2 => n238, B => 
                           valid_data_port, C => write_en, Y => n235);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_0_port, A2 => n17, B1 => 
                           data_in(0), B2 => n29, Y => n234);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_1_port, A2 => n17, B1 => 
                           data_in(1), B2 => n29, Y => n233);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_2_port, A2 => n17, B1 => 
                           data_in(2), B2 => n29, Y => n232);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_3_port, A2 => n17, B1 => 
                           data_in(3), B2 => n29, Y => n231);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_4_port, A2 => n17, B1 => 
                           data_in(4), B2 => n27, Y => n230);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_5_port, A2 => n17, B1 => 
                           data_in(5), B2 => n27, Y => n229);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_6_port, A2 => n17, B1 => 
                           data_in(6), B2 => n27, Y => n228);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_7_port, A2 => n17, B1 => 
                           data_in(7), B2 => n27, Y => n227);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_8_port, A2 => n17, B1 => 
                           data_in(8), B2 => n27, Y => n226);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_9_port, A2 => n17, B1 => 
                           data_in(9), B2 => n27, Y => n225);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_10_port, A2 => n17, B1 => 
                           data_in(10), B2 => n27, Y => n224);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_11_port, A2 => n17, B1 => 
                           data_in(11), B2 => n27, Y => n223);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_12_port, A2 => n17, B1 => 
                           data_in(12), B2 => n27, Y => n222);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_13_port, A2 => n17, B1 => 
                           data_in(13), B2 => n27, Y => n221);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_14_port, A2 => n17, B1 => 
                           data_in(14), B2 => n27, Y => n220);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_15_port, A2 => n17, B1 => 
                           data_in(15), B2 => n27, Y => n219);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_16_port, A2 => n17, B1 => 
                           data_in(16), B2 => n25, Y => n218);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_17_port, A2 => n17, B1 => 
                           data_in(17), B2 => n25, Y => n217);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_18_port, A2 => n17, B1 => 
                           data_in(18), B2 => n25, Y => n216);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_19_port, A2 => n17, B1 => 
                           data_in(19), B2 => n25, Y => n215);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_20_port, A2 => n17, B1 => 
                           data_in(20), B2 => n25, Y => n214);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_21_port, A2 => n17, B1 => 
                           data_in(21), B2 => n25, Y => n213);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_22_port, A2 => n17, B1 => 
                           data_in(22), B2 => n25, Y => n212);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_23_port, A2 => n17, B1 => 
                           data_in(23), B2 => n25, Y => n211);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_24_port, A2 => n17, B1 => 
                           data_in(24), B2 => n25, Y => n210);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_25_port, A2 => n17, B1 => 
                           data_in(25), B2 => n25, Y => n209);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_26_port, A2 => n17, B1 => 
                           data_in(26), B2 => n25, Y => n208);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_27_port, A2 => n17, B1 => 
                           data_in(27), B2 => n25, Y => n207);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_28_port, A2 => n17, B1 => 
                           data_in(28), B2 => n23, Y => n206);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_29_port, A2 => n17, B1 => 
                           data_in(29), B2 => n23, Y => n205);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_30_port, A2 => n17, B1 => 
                           data_in(30), B2 => n23, Y => n204);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_31_port, A2 => n17, B1 => 
                           data_in(31), B2 => n23, Y => n203);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_32_port, A2 => n17, B1 => 
                           data_in(32), B2 => n23, Y => n202);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_33_port, A2 => n17, B1 => 
                           data_in(33), B2 => n23, Y => n201);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_34_port, A2 => n17, B1 => 
                           data_in(34), B2 => n23, Y => n200);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_35_port, A2 => n17, B1 => 
                           data_in(35), B2 => n23, Y => n199);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_36_port, A2 => n17, B1 => 
                           data_in(36), B2 => n23, Y => n198);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_37_port, A2 => n17, B1 => 
                           data_in(37), B2 => n23, Y => n197);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_38_port, A2 => n17, B1 => 
                           data_in(38), B2 => n23, Y => n196);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_39_port, A2 => n17, B1 => 
                           data_in(39), B2 => n23, Y => n195);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_40_port, A2 => n17, B1 => 
                           data_in(40), B2 => n21, Y => n194);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_41_port, A2 => n17, B1 => 
                           data_in(41), B2 => n21, Y => n193);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_42_port, A2 => n17, B1 => 
                           data_in(42), B2 => n21, Y => n192);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_43_port, A2 => n17, B1 => 
                           data_in(43), B2 => n21, Y => n191);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_44_port, A2 => n17, B1 => 
                           data_in(44), B2 => n21, Y => n190);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_45_port, A2 => n17, B1 => 
                           data_in(45), B2 => n21, Y => n189);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_46_port, A2 => n17, B1 => 
                           data_in(46), B2 => n21, Y => n188);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_47_port, A2 => n17, B1 => 
                           data_in(47), B2 => n21, Y => n187);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_48_port, A2 => n17, B1 => 
                           data_in(48), B2 => n21, Y => n186);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_49_port, A2 => n17, B1 => 
                           data_in(49), B2 => n21, Y => n185);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_50_port, A2 => n17, B1 => 
                           data_in(50), B2 => n21, Y => n184);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_51_port, A2 => n17, B1 => 
                           data_in(51), B2 => n21, Y => n183);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_52_port, A2 => n17, B1 => 
                           data_in(52), B2 => n19, Y => n182);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_53_port, A2 => n17, B1 => 
                           data_in(53), B2 => n19, Y => n181);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_54_port, A2 => n17, B1 => 
                           data_in(54), B2 => n19, Y => n180);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_55_port, A2 => n17, B1 => 
                           data_in(55), B2 => n19, Y => n179);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_56_port, A2 => n17, B1 => 
                           data_in(56), B2 => n19, Y => n178);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_57_port, A2 => n17, B1 => 
                           data_in(57), B2 => n19, Y => n177);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_58_port, A2 => n17, B1 => 
                           data_in(58), B2 => n19, Y => n176);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_59_port, A2 => n17, B1 => 
                           data_in(59), B2 => n19, Y => n175);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_60_port, A2 => n17, B1 => 
                           data_in(60), B2 => n19, Y => n174);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_61_port, A2 => n17, B1 => 
                           data_in(61), B2 => n19, Y => n173);
   U67 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_62_port, A2 => n17, B1 => 
                           data_in(62), B2 => n19, Y => n172);
   U68 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_63_port, A2 => n17, B1 => 
                           data_in(63), B2 => n19, Y => n171);
   U70 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N9, Y => n237);
   U71 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_0_port, A2 => n3, B1 => 
                           data_in(0), B2 => n15, Y => n170);
   U72 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_1_port, A2 => n3, B1 => 
                           data_in(1), B2 => n15, Y => n169);
   U73 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_2_port, A2 => n3, B1 => 
                           data_in(2), B2 => n15, Y => n168);
   U74 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_3_port, A2 => n3, B1 => 
                           data_in(3), B2 => n15, Y => n167);
   U75 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_4_port, A2 => n3, B1 => 
                           data_in(4), B2 => n13, Y => n166);
   U76 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_5_port, A2 => n3, B1 => 
                           data_in(5), B2 => n13, Y => n165);
   U77 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_6_port, A2 => n3, B1 => 
                           data_in(6), B2 => n13, Y => n164);
   U78 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_7_port, A2 => n3, B1 => 
                           data_in(7), B2 => n13, Y => n163);
   U79 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_8_port, A2 => n3, B1 => 
                           data_in(8), B2 => n13, Y => n162);
   U80 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_9_port, A2 => n3, B1 => 
                           data_in(9), B2 => n13, Y => n161);
   U81 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_10_port, A2 => n3, B1 => 
                           data_in(10), B2 => n13, Y => n160);
   U82 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_11_port, A2 => n3, B1 => 
                           data_in(11), B2 => n13, Y => n159);
   U83 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_12_port, A2 => n3, B1 => 
                           data_in(12), B2 => n13, Y => n157);
   U84 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_13_port, A2 => n3, B1 => 
                           data_in(13), B2 => n13, Y => n155);
   U85 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_14_port, A2 => n3, B1 => 
                           data_in(14), B2 => n13, Y => n153);
   U86 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_15_port, A2 => n3, B1 => 
                           data_in(15), B2 => n13, Y => n151);
   U87 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_16_port, A2 => n3, B1 => 
                           data_in(16), B2 => n11, Y => n149);
   U88 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_17_port, A2 => n3, B1 => 
                           data_in(17), B2 => n11, Y => n147);
   U89 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_18_port, A2 => n3, B1 => 
                           data_in(18), B2 => n11, Y => n145);
   U90 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_19_port, A2 => n3, B1 => 
                           data_in(19), B2 => n11, Y => n143);
   U91 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_20_port, A2 => n3, B1 => 
                           data_in(20), B2 => n11, Y => n141);
   U92 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_21_port, A2 => n3, B1 => 
                           data_in(21), B2 => n11, Y => n139);
   U93 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_22_port, A2 => n3, B1 => 
                           data_in(22), B2 => n11, Y => n137);
   U94 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_23_port, A2 => n3, B1 => 
                           data_in(23), B2 => n11, Y => n135);
   U95 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_24_port, A2 => n3, B1 => 
                           data_in(24), B2 => n11, Y => n133);
   U96 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_25_port, A2 => n3, B1 => 
                           data_in(25), B2 => n11, Y => n131);
   U97 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_26_port, A2 => n3, B1 => 
                           data_in(26), B2 => n11, Y => n129);
   U98 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_27_port, A2 => n3, B1 => 
                           data_in(27), B2 => n11, Y => n127);
   U99 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_28_port, A2 => n3, B1 => 
                           data_in(28), B2 => n9_port, Y => n125);
   U100 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_29_port, A2 => n3, B1 => 
                           data_in(29), B2 => n9_port, Y => n123);
   U101 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_30_port, A2 => n3, B1 => 
                           data_in(30), B2 => n9_port, Y => n121);
   U102 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_31_port, A2 => n3, B1 => 
                           data_in(31), B2 => n9_port, Y => n119);
   U103 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_32_port, A2 => n3, B1 => 
                           data_in(32), B2 => n9_port, Y => n117);
   U104 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_33_port, A2 => n3, B1 => 
                           data_in(33), B2 => n9_port, Y => n115);
   U105 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_34_port, A2 => n3, B1 => 
                           data_in(34), B2 => n9_port, Y => n113);
   U106 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_35_port, A2 => n3, B1 => 
                           data_in(35), B2 => n9_port, Y => n111);
   U107 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_36_port, A2 => n3, B1 => 
                           data_in(36), B2 => n9_port, Y => n109);
   U108 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_37_port, A2 => n3, B1 => 
                           data_in(37), B2 => n9_port, Y => n107);
   U109 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_38_port, A2 => n3, B1 => 
                           data_in(38), B2 => n9_port, Y => n105);
   U110 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_39_port, A2 => n3, B1 => 
                           data_in(39), B2 => n9_port, Y => n103);
   U111 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_40_port, A2 => n3, B1 => 
                           data_in(40), B2 => n7_port, Y => n101);
   U112 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_41_port, A2 => n3, B1 => 
                           data_in(41), B2 => n7_port, Y => n99);
   U113 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_42_port, A2 => n3, B1 => 
                           data_in(42), B2 => n7_port, Y => n97);
   U114 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_43_port, A2 => n3, B1 => 
                           data_in(43), B2 => n7_port, Y => n95);
   U115 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_44_port, A2 => n3, B1 => 
                           data_in(44), B2 => n7_port, Y => n93);
   U116 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_45_port, A2 => n3, B1 => 
                           data_in(45), B2 => n7_port, Y => n91);
   U117 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_46_port, A2 => n3, B1 => 
                           data_in(46), B2 => n7_port, Y => n89);
   U118 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_47_port, A2 => n3, B1 => 
                           data_in(47), B2 => n7_port, Y => n87);
   U119 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_48_port, A2 => n3, B1 => 
                           data_in(48), B2 => n7_port, Y => n85);
   U120 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_49_port, A2 => n3, B1 => 
                           data_in(49), B2 => n7_port, Y => n83);
   U121 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_50_port, A2 => n3, B1 => 
                           data_in(50), B2 => n7_port, Y => n81);
   U122 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_51_port, A2 => n3, B1 => 
                           data_in(51), B2 => n7_port, Y => n79);
   U123 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_52_port, A2 => n3, B1 => 
                           data_in(52), B2 => n5, Y => n77);
   U124 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_53_port, A2 => n3, B1 => 
                           data_in(53), B2 => n5, Y => n75);
   U125 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_54_port, A2 => n3, B1 => 
                           data_in(54), B2 => n5, Y => n73);
   U126 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_55_port, A2 => n3, B1 => 
                           data_in(55), B2 => n5, Y => n71);
   U127 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_56_port, A2 => n3, B1 => 
                           data_in(56), B2 => n5, Y => n69);
   U128 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_57_port, A2 => n3, B1 => 
                           data_in(57), B2 => n5, Y => n67);
   U129 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_58_port, A2 => n3, B1 => 
                           data_in(58), B2 => n5, Y => n65);
   U130 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_59_port, A2 => n3, B1 => 
                           data_in(59), B2 => n5, Y => n63);
   U131 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_60_port, A2 => n3, B1 => 
                           data_in(60), B2 => n5, Y => n61);
   U132 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_61_port, A2 => n3, B1 => 
                           data_in(61), B2 => n5, Y => n59);
   U133 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_62_port, A2 => n3, B1 => 
                           data_in(62), B2 => n5, Y => n57);
   U134 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_63_port, A2 => n3, B1 => 
                           data_in(63), B2 => n5, Y => n55);
   U136 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N7, Y => n236);
   U137 : OAI22xp5_ASAP7_75t_R port map( A1 => n31, A2 => read_en, B1 => n43, 
                           B2 => n47, Y => n53);
   U139 : OAI22xp5_ASAP7_75t_R port map( A1 => N9, A2 => n49, B1 => write_en, 
                           B2 => N7, Y => n51);
   write_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK 
                           => clk, RESET => n45, SET => n1, QN => N7);
   fifo_reg_1_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n55, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_63_port);
   fifo_reg_1_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n57, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_62_port);
   fifo_reg_1_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n59, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_61_port);
   fifo_reg_1_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n61, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_60_port);
   fifo_reg_0_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n171, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_63_port);
   fifo_reg_0_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n172, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_62_port);
   fifo_reg_0_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n173, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_61_port);
   fifo_reg_0_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n174, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_60_port);
   fifo_reg_1_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n167, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_3_port);
   fifo_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n168, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_2_port);
   fifo_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n169, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_1_port);
   fifo_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n170, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_0_port);
   fifo_reg_1_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n63, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_59_port);
   fifo_reg_1_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n65, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_58_port);
   fifo_reg_1_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n67, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_57_port);
   fifo_reg_1_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n69, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_56_port);
   fifo_reg_1_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n71, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_55_port);
   fifo_reg_1_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n73, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_54_port);
   fifo_reg_1_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n75, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_53_port);
   fifo_reg_1_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n77, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_52_port);
   fifo_reg_1_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_51_port);
   fifo_reg_1_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_50_port);
   fifo_reg_1_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_49_port);
   fifo_reg_1_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_48_port);
   fifo_reg_1_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_47_port);
   fifo_reg_1_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_46_port);
   fifo_reg_1_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_45_port);
   fifo_reg_1_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_44_port);
   fifo_reg_1_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_43_port);
   fifo_reg_1_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_42_port);
   fifo_reg_1_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_41_port);
   fifo_reg_1_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_40_port);
   fifo_reg_1_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_39_port);
   fifo_reg_1_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_38_port);
   fifo_reg_1_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_37_port);
   fifo_reg_1_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_36_port);
   fifo_reg_1_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_35_port);
   fifo_reg_1_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_34_port);
   fifo_reg_1_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n115, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_33_port);
   fifo_reg_1_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n117, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_32_port);
   fifo_reg_1_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n119, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_31_port);
   fifo_reg_1_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n121, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_30_port);
   fifo_reg_1_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n123, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_29_port);
   fifo_reg_1_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n125, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_28_port);
   fifo_reg_1_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n127, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_27_port);
   fifo_reg_1_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n129, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_26_port);
   fifo_reg_1_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n131, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_25_port);
   fifo_reg_1_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n133, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_24_port);
   fifo_reg_1_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n135, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_23_port);
   fifo_reg_1_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n137, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_22_port);
   fifo_reg_1_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n139, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_21_port);
   fifo_reg_1_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n141, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_20_port);
   fifo_reg_1_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n143, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_19_port);
   fifo_reg_1_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n145, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_18_port);
   fifo_reg_1_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n147, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_17_port);
   fifo_reg_1_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n149, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_16_port);
   fifo_reg_1_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n151, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_15_port);
   fifo_reg_1_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n153, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_14_port);
   fifo_reg_1_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n155, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_13_port);
   fifo_reg_1_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n157, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_12_port);
   fifo_reg_1_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n159, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_11_port);
   fifo_reg_1_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n160, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_10_port);
   fifo_reg_1_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n161, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_9_port);
   fifo_reg_1_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n162, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_8_port);
   fifo_reg_1_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n163, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_7_port);
   fifo_reg_1_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n164, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_6_port);
   fifo_reg_1_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n165, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_5_port);
   fifo_reg_1_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n166, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_4_port);
   fifo_reg_0_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n231, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_3_port);
   fifo_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n232, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_2_port);
   fifo_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n233, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_1_port);
   fifo_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n234, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_0_port);
   fifo_reg_0_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n175, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_59_port);
   fifo_reg_0_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n176, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_58_port);
   fifo_reg_0_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n177, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_57_port);
   fifo_reg_0_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n178, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_56_port);
   fifo_reg_0_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n179, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_55_port);
   fifo_reg_0_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n180, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_54_port);
   fifo_reg_0_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n181, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_53_port);
   fifo_reg_0_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n182, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_52_port);
   fifo_reg_0_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n183, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_51_port);
   fifo_reg_0_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n184, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_50_port);
   fifo_reg_0_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n185, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_49_port);
   fifo_reg_0_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n186, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_48_port);
   fifo_reg_0_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n187, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_47_port);
   fifo_reg_0_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n188, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_46_port);
   fifo_reg_0_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n189, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_45_port);
   fifo_reg_0_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n190, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_44_port);
   fifo_reg_0_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n191, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_43_port);
   fifo_reg_0_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n192, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_42_port);
   fifo_reg_0_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n193, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_41_port);
   fifo_reg_0_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n194, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_40_port);
   fifo_reg_0_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n195, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_39_port);
   fifo_reg_0_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n196, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_38_port);
   fifo_reg_0_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n197, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_37_port);
   fifo_reg_0_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n198, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_36_port);
   fifo_reg_0_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n199, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_35_port);
   fifo_reg_0_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n200, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_34_port);
   fifo_reg_0_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n201, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_33_port);
   fifo_reg_0_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n202, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_32_port);
   fifo_reg_0_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n203, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_31_port);
   fifo_reg_0_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n204, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_30_port);
   fifo_reg_0_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n205, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_29_port);
   fifo_reg_0_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n206, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_28_port);
   fifo_reg_0_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n207, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_27_port);
   fifo_reg_0_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n208, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_26_port);
   fifo_reg_0_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n209, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_25_port);
   fifo_reg_0_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n210, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_24_port);
   fifo_reg_0_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n211, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_23_port);
   fifo_reg_0_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n212, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_22_port);
   fifo_reg_0_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n213, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_21_port);
   fifo_reg_0_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n214, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_20_port);
   fifo_reg_0_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n215, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_19_port);
   fifo_reg_0_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n216, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_18_port);
   fifo_reg_0_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n217, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_17_port);
   fifo_reg_0_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n218, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_16_port);
   fifo_reg_0_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n219, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_15_port);
   fifo_reg_0_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n220, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_14_port);
   fifo_reg_0_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n221, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_13_port);
   fifo_reg_0_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n222, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_12_port);
   fifo_reg_0_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n223, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_11_port);
   fifo_reg_0_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n224, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_10_port);
   fifo_reg_0_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n225, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_9_port);
   fifo_reg_0_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n226, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_8_port);
   fifo_reg_0_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n227, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_7_port);
   fifo_reg_0_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n228, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_6_port);
   fifo_reg_0_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n229, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_5_port);
   fifo_reg_0_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n230, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_4_port);
   read_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK 
                           => clk, RESET => n45, SET => n1, QN => 
                           read_pointer_0_port);
   valid_data_reg : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n235, CLK => clk, 
                           RESET => n45, SET => n1, QN => valid_data_port);
   U69 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U135 : INVx3_ASAP7_75t_R port map( A => rst, Y => n45);
   U138 : INVx1_ASAP7_75t_R port map( A => n29, Y => n17);
   U140 : INVx1_ASAP7_75t_R port map( A => n15, Y => n3);
   U141 : INVx1_ASAP7_75t_R port map( A => n31, Y => n43);
   U142 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n29);
   U207 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n15);
   U208 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n27);
   U209 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n25);
   U210 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n23);
   U211 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n21);
   U212 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n19);
   U213 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n13);
   U214 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n11);
   U215 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n9_port);
   U216 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n7_port);
   U217 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n5);
   U218 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n31);
   U219 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n33);
   U220 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n41);
   U221 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n39);
   U222 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n37);
   U223 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n35);
   U224 : INVx1_ASAP7_75t_R port map( A => read_en, Y => n47);
   U225 : INVx1_ASAP7_75t_R port map( A => N7, Y => N9);
   U226 : INVx1_ASAP7_75t_R port map( A => write_en, Y => n49);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity fifo_buff_depth2_3 is

   port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, clk, 
         rst : in std_logic;  data_out : out std_logic_vector (63 downto 0);  
         valid_data : out std_logic);

end fifo_buff_depth2_3;

architecture SYN_rtl of fifo_buff_depth2_3 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx3_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal valid_data_port, read_pointer_0_port, fifo_1_63_port, fifo_1_62_port,
      fifo_1_61_port, fifo_1_60_port, fifo_1_59_port, fifo_1_58_port, 
      fifo_1_57_port, fifo_1_56_port, fifo_1_55_port, fifo_1_54_port, 
      fifo_1_53_port, fifo_1_52_port, fifo_1_51_port, fifo_1_50_port, 
      fifo_1_49_port, fifo_1_48_port, fifo_1_47_port, fifo_1_46_port, 
      fifo_1_45_port, fifo_1_44_port, fifo_1_43_port, fifo_1_42_port, 
      fifo_1_41_port, fifo_1_40_port, fifo_1_39_port, fifo_1_38_port, 
      fifo_1_37_port, fifo_1_36_port, fifo_1_35_port, fifo_1_34_port, 
      fifo_1_33_port, fifo_1_32_port, fifo_1_31_port, fifo_1_30_port, 
      fifo_1_29_port, fifo_1_28_port, fifo_1_27_port, fifo_1_26_port, 
      fifo_1_25_port, fifo_1_24_port, fifo_1_23_port, fifo_1_22_port, 
      fifo_1_21_port, fifo_1_20_port, fifo_1_19_port, fifo_1_18_port, 
      fifo_1_17_port, fifo_1_16_port, fifo_1_15_port, fifo_1_14_port, 
      fifo_1_13_port, fifo_1_12_port, fifo_1_11_port, fifo_1_10_port, 
      fifo_1_9_port, fifo_1_8_port, fifo_1_7_port, fifo_1_6_port, fifo_1_5_port
      , fifo_1_4_port, fifo_1_3_port, fifo_1_2_port, fifo_1_1_port, 
      fifo_1_0_port, fifo_0_63_port, fifo_0_62_port, fifo_0_61_port, 
      fifo_0_60_port, fifo_0_59_port, fifo_0_58_port, fifo_0_57_port, 
      fifo_0_56_port, fifo_0_55_port, fifo_0_54_port, fifo_0_53_port, 
      fifo_0_52_port, fifo_0_51_port, fifo_0_50_port, fifo_0_49_port, 
      fifo_0_48_port, fifo_0_47_port, fifo_0_46_port, fifo_0_45_port, 
      fifo_0_44_port, fifo_0_43_port, fifo_0_42_port, fifo_0_41_port, 
      fifo_0_40_port, fifo_0_39_port, fifo_0_38_port, fifo_0_37_port, 
      fifo_0_36_port, fifo_0_35_port, fifo_0_34_port, fifo_0_33_port, 
      fifo_0_32_port, fifo_0_31_port, fifo_0_30_port, fifo_0_29_port, 
      fifo_0_28_port, fifo_0_27_port, fifo_0_26_port, fifo_0_25_port, 
      fifo_0_24_port, fifo_0_23_port, fifo_0_22_port, fifo_0_21_port, 
      fifo_0_20_port, fifo_0_19_port, fifo_0_18_port, fifo_0_17_port, 
      fifo_0_16_port, fifo_0_15_port, fifo_0_14_port, fifo_0_13_port, 
      fifo_0_12_port, fifo_0_11_port, fifo_0_10_port, fifo_0_9_port, 
      fifo_0_8_port, fifo_0_7_port, fifo_0_6_port, fifo_0_5_port, fifo_0_4_port
      , fifo_0_3_port, fifo_0_2_port, fifo_0_1_port, fifo_0_0_port, N7, N9, n1,
      n3, n5, n7_port, n9_port, n11, n13, n15, n17, n19, n21, n23, n25, n27, 
      n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57
      , n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, 
      n87, n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, n111, 
      n113, n115, n117, n119, n121, n123, n125, n127, n129, n131, n133, n135, 
      n137, n139, n141, n143, n145, n147, n149, n151, n153, n155, n157, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238 : std_logic;

begin
   valid_data <= valid_data_port;
   
   U4 : XOR2xp5_ASAP7_75t_R port map( A => N7, B => n43, Y => n238);
   U143 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_9_port, B1 => 
                           n43, B2 => fifo_0_9_port, Y => data_out(9));
   U144 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_8_port, B1 => 
                           n43, B2 => fifo_0_8_port, Y => data_out(8));
   U145 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_7_port, B1 => 
                           n43, B2 => fifo_0_7_port, Y => data_out(7));
   U146 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_6_port, B1 => 
                           n43, B2 => fifo_0_6_port, Y => data_out(6));
   U147 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_63_port, B1 => 
                           n43, B2 => fifo_0_63_port, Y => data_out(63));
   U148 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_62_port, B1 => 
                           n43, B2 => fifo_0_62_port, Y => data_out(62));
   U149 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_61_port, B1 => 
                           n43, B2 => fifo_0_61_port, Y => data_out(61));
   U150 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_60_port, B1 => 
                           n43, B2 => fifo_0_60_port, Y => data_out(60));
   U151 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_5_port, B1 => 
                           n43, B2 => fifo_0_5_port, Y => data_out(5));
   U152 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_59_port, B1 => 
                           n43, B2 => fifo_0_59_port, Y => data_out(59));
   U153 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_58_port, B1 => 
                           n43, B2 => fifo_0_58_port, Y => data_out(58));
   U154 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_57_port, B1 => 
                           n43, B2 => fifo_0_57_port, Y => data_out(57));
   U155 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_56_port, B1 => 
                           n43, B2 => fifo_0_56_port, Y => data_out(56));
   U156 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_55_port, B1 => 
                           n43, B2 => fifo_0_55_port, Y => data_out(55));
   U157 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_54_port, B1 => 
                           n43, B2 => fifo_0_54_port, Y => data_out(54));
   U158 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_53_port, B1 => 
                           n43, B2 => fifo_0_53_port, Y => data_out(53));
   U159 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_52_port, B1 => 
                           n43, B2 => fifo_0_52_port, Y => data_out(52));
   U160 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_51_port, B1 => 
                           n43, B2 => fifo_0_51_port, Y => data_out(51));
   U161 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_50_port, B1 => 
                           n43, B2 => fifo_0_50_port, Y => data_out(50));
   U162 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_4_port, B1 => 
                           n43, B2 => fifo_0_4_port, Y => data_out(4));
   U163 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_49_port, B1 => 
                           n43, B2 => fifo_0_49_port, Y => data_out(49));
   U164 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_48_port, B1 => 
                           n43, B2 => fifo_0_48_port, Y => data_out(48));
   U165 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_47_port, B1 => 
                           n43, B2 => fifo_0_47_port, Y => data_out(47));
   U166 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_46_port, B1 => 
                           n43, B2 => fifo_0_46_port, Y => data_out(46));
   U167 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_45_port, B1 => 
                           n43, B2 => fifo_0_45_port, Y => data_out(45));
   U168 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_44_port, B1 => 
                           n43, B2 => fifo_0_44_port, Y => data_out(44));
   U169 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_43_port, B1 => 
                           n43, B2 => fifo_0_43_port, Y => data_out(43));
   U170 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_42_port, B1 => 
                           n43, B2 => fifo_0_42_port, Y => data_out(42));
   U171 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_41_port, B1 => 
                           n43, B2 => fifo_0_41_port, Y => data_out(41));
   U172 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_40_port, B1 => 
                           n43, B2 => fifo_0_40_port, Y => data_out(40));
   U173 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_3_port, B1 => 
                           n43, B2 => fifo_0_3_port, Y => data_out(3));
   U174 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_39_port, B1 => 
                           n43, B2 => fifo_0_39_port, Y => data_out(39));
   U175 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_38_port, B1 => 
                           n43, B2 => fifo_0_38_port, Y => data_out(38));
   U176 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_37_port, B1 => 
                           n43, B2 => fifo_0_37_port, Y => data_out(37));
   U177 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_36_port, B1 => 
                           n43, B2 => fifo_0_36_port, Y => data_out(36));
   U178 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_35_port, B1 => 
                           n43, B2 => fifo_0_35_port, Y => data_out(35));
   U179 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_34_port, B1 => 
                           n43, B2 => fifo_0_34_port, Y => data_out(34));
   U180 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_33_port, B1 => 
                           n43, B2 => fifo_0_33_port, Y => data_out(33));
   U181 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_32_port, B1 => 
                           n43, B2 => fifo_0_32_port, Y => data_out(32));
   U182 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_31_port, B1 => 
                           n43, B2 => fifo_0_31_port, Y => data_out(31));
   U183 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_30_port, B1 => 
                           n43, B2 => fifo_0_30_port, Y => data_out(30));
   U184 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_2_port, B1 => 
                           n43, B2 => fifo_0_2_port, Y => data_out(2));
   U185 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_29_port, B1 => 
                           n43, B2 => fifo_0_29_port, Y => data_out(29));
   U186 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_28_port, B1 => 
                           n43, B2 => fifo_0_28_port, Y => data_out(28));
   U187 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_27_port, B1 => 
                           n43, B2 => fifo_0_27_port, Y => data_out(27));
   U188 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_26_port, B1 => 
                           n43, B2 => fifo_0_26_port, Y => data_out(26));
   U189 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_25_port, B1 => 
                           n43, B2 => fifo_0_25_port, Y => data_out(25));
   U190 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_24_port, B1 => 
                           n43, B2 => fifo_0_24_port, Y => data_out(24));
   U191 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_23_port, B1 => 
                           n43, B2 => fifo_0_23_port, Y => data_out(23));
   U192 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_22_port, B1 => 
                           n43, B2 => fifo_0_22_port, Y => data_out(22));
   U193 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_21_port, B1 => 
                           n43, B2 => fifo_0_21_port, Y => data_out(21));
   U194 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_20_port, B1 => 
                           n43, B2 => fifo_0_20_port, Y => data_out(20));
   U195 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_1_port, B1 => 
                           n43, B2 => fifo_0_1_port, Y => data_out(1));
   U196 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_19_port, B1 => 
                           n43, B2 => fifo_0_19_port, Y => data_out(19));
   U197 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_18_port, B1 => 
                           n43, B2 => fifo_0_18_port, Y => data_out(18));
   U198 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_17_port, B1 => 
                           n43, B2 => fifo_0_17_port, Y => data_out(17));
   U199 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_16_port, B1 => 
                           n43, B2 => fifo_0_16_port, Y => data_out(16));
   U200 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_15_port, B1 => 
                           n43, B2 => fifo_0_15_port, Y => data_out(15));
   U201 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_14_port, B1 => 
                           n43, B2 => fifo_0_14_port, Y => data_out(14));
   U202 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_13_port, B1 => 
                           n43, B2 => fifo_0_13_port, Y => data_out(13));
   U203 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_12_port, B1 => 
                           n43, B2 => fifo_0_12_port, Y => data_out(12));
   U204 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_11_port, B1 => 
                           n43, B2 => fifo_0_11_port, Y => data_out(11));
   U205 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_10_port, B1 => 
                           n43, B2 => fifo_0_10_port, Y => data_out(10));
   U206 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_0_port, B1 => 
                           n43, B2 => fifo_0_0_port, Y => data_out(0));
   U3 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n45, A2 => n238, B => 
                           valid_data_port, C => write_en, Y => n235);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_0_port, A2 => n17, B1 => 
                           data_in(0), B2 => n29, Y => n234);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_1_port, A2 => n17, B1 => 
                           data_in(1), B2 => n29, Y => n233);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_2_port, A2 => n17, B1 => 
                           data_in(2), B2 => n29, Y => n232);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_3_port, A2 => n17, B1 => 
                           data_in(3), B2 => n29, Y => n231);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_4_port, A2 => n17, B1 => 
                           data_in(4), B2 => n27, Y => n230);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_5_port, A2 => n17, B1 => 
                           data_in(5), B2 => n27, Y => n229);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_6_port, A2 => n17, B1 => 
                           data_in(6), B2 => n27, Y => n228);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_7_port, A2 => n17, B1 => 
                           data_in(7), B2 => n27, Y => n227);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_8_port, A2 => n17, B1 => 
                           data_in(8), B2 => n27, Y => n226);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_9_port, A2 => n17, B1 => 
                           data_in(9), B2 => n27, Y => n225);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_10_port, A2 => n17, B1 => 
                           data_in(10), B2 => n27, Y => n224);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_11_port, A2 => n17, B1 => 
                           data_in(11), B2 => n27, Y => n223);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_12_port, A2 => n17, B1 => 
                           data_in(12), B2 => n27, Y => n222);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_13_port, A2 => n17, B1 => 
                           data_in(13), B2 => n27, Y => n221);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_14_port, A2 => n17, B1 => 
                           data_in(14), B2 => n27, Y => n220);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_15_port, A2 => n17, B1 => 
                           data_in(15), B2 => n27, Y => n219);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_16_port, A2 => n17, B1 => 
                           data_in(16), B2 => n25, Y => n218);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_17_port, A2 => n17, B1 => 
                           data_in(17), B2 => n25, Y => n217);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_18_port, A2 => n17, B1 => 
                           data_in(18), B2 => n25, Y => n216);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_19_port, A2 => n17, B1 => 
                           data_in(19), B2 => n25, Y => n215);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_20_port, A2 => n17, B1 => 
                           data_in(20), B2 => n25, Y => n214);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_21_port, A2 => n17, B1 => 
                           data_in(21), B2 => n25, Y => n213);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_22_port, A2 => n17, B1 => 
                           data_in(22), B2 => n25, Y => n212);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_23_port, A2 => n17, B1 => 
                           data_in(23), B2 => n25, Y => n211);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_24_port, A2 => n17, B1 => 
                           data_in(24), B2 => n25, Y => n210);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_25_port, A2 => n17, B1 => 
                           data_in(25), B2 => n25, Y => n209);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_26_port, A2 => n17, B1 => 
                           data_in(26), B2 => n25, Y => n208);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_27_port, A2 => n17, B1 => 
                           data_in(27), B2 => n25, Y => n207);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_28_port, A2 => n17, B1 => 
                           data_in(28), B2 => n23, Y => n206);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_29_port, A2 => n17, B1 => 
                           data_in(29), B2 => n23, Y => n205);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_30_port, A2 => n17, B1 => 
                           data_in(30), B2 => n23, Y => n204);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_31_port, A2 => n17, B1 => 
                           data_in(31), B2 => n23, Y => n203);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_32_port, A2 => n17, B1 => 
                           data_in(32), B2 => n23, Y => n202);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_33_port, A2 => n17, B1 => 
                           data_in(33), B2 => n23, Y => n201);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_34_port, A2 => n17, B1 => 
                           data_in(34), B2 => n23, Y => n200);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_35_port, A2 => n17, B1 => 
                           data_in(35), B2 => n23, Y => n199);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_36_port, A2 => n17, B1 => 
                           data_in(36), B2 => n23, Y => n198);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_37_port, A2 => n17, B1 => 
                           data_in(37), B2 => n23, Y => n197);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_38_port, A2 => n17, B1 => 
                           data_in(38), B2 => n23, Y => n196);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_39_port, A2 => n17, B1 => 
                           data_in(39), B2 => n23, Y => n195);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_40_port, A2 => n17, B1 => 
                           data_in(40), B2 => n21, Y => n194);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_41_port, A2 => n17, B1 => 
                           data_in(41), B2 => n21, Y => n193);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_42_port, A2 => n17, B1 => 
                           data_in(42), B2 => n21, Y => n192);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_43_port, A2 => n17, B1 => 
                           data_in(43), B2 => n21, Y => n191);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_44_port, A2 => n17, B1 => 
                           data_in(44), B2 => n21, Y => n190);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_45_port, A2 => n17, B1 => 
                           data_in(45), B2 => n21, Y => n189);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_46_port, A2 => n17, B1 => 
                           data_in(46), B2 => n21, Y => n188);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_47_port, A2 => n17, B1 => 
                           data_in(47), B2 => n21, Y => n187);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_48_port, A2 => n17, B1 => 
                           data_in(48), B2 => n21, Y => n186);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_49_port, A2 => n17, B1 => 
                           data_in(49), B2 => n21, Y => n185);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_50_port, A2 => n17, B1 => 
                           data_in(50), B2 => n21, Y => n184);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_51_port, A2 => n17, B1 => 
                           data_in(51), B2 => n21, Y => n183);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_52_port, A2 => n17, B1 => 
                           data_in(52), B2 => n19, Y => n182);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_53_port, A2 => n17, B1 => 
                           data_in(53), B2 => n19, Y => n181);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_54_port, A2 => n17, B1 => 
                           data_in(54), B2 => n19, Y => n180);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_55_port, A2 => n17, B1 => 
                           data_in(55), B2 => n19, Y => n179);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_56_port, A2 => n17, B1 => 
                           data_in(56), B2 => n19, Y => n178);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_57_port, A2 => n17, B1 => 
                           data_in(57), B2 => n19, Y => n177);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_58_port, A2 => n17, B1 => 
                           data_in(58), B2 => n19, Y => n176);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_59_port, A2 => n17, B1 => 
                           data_in(59), B2 => n19, Y => n175);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_60_port, A2 => n17, B1 => 
                           data_in(60), B2 => n19, Y => n174);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_61_port, A2 => n17, B1 => 
                           data_in(61), B2 => n19, Y => n173);
   U67 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_62_port, A2 => n17, B1 => 
                           data_in(62), B2 => n19, Y => n172);
   U68 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_63_port, A2 => n17, B1 => 
                           data_in(63), B2 => n19, Y => n171);
   U70 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N9, Y => n237);
   U71 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_0_port, A2 => n3, B1 => 
                           data_in(0), B2 => n15, Y => n170);
   U72 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_1_port, A2 => n3, B1 => 
                           data_in(1), B2 => n15, Y => n169);
   U73 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_2_port, A2 => n3, B1 => 
                           data_in(2), B2 => n15, Y => n168);
   U74 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_3_port, A2 => n3, B1 => 
                           data_in(3), B2 => n15, Y => n167);
   U75 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_4_port, A2 => n3, B1 => 
                           data_in(4), B2 => n13, Y => n166);
   U76 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_5_port, A2 => n3, B1 => 
                           data_in(5), B2 => n13, Y => n165);
   U77 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_6_port, A2 => n3, B1 => 
                           data_in(6), B2 => n13, Y => n164);
   U78 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_7_port, A2 => n3, B1 => 
                           data_in(7), B2 => n13, Y => n163);
   U79 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_8_port, A2 => n3, B1 => 
                           data_in(8), B2 => n13, Y => n162);
   U80 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_9_port, A2 => n3, B1 => 
                           data_in(9), B2 => n13, Y => n161);
   U81 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_10_port, A2 => n3, B1 => 
                           data_in(10), B2 => n13, Y => n160);
   U82 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_11_port, A2 => n3, B1 => 
                           data_in(11), B2 => n13, Y => n159);
   U83 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_12_port, A2 => n3, B1 => 
                           data_in(12), B2 => n13, Y => n157);
   U84 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_13_port, A2 => n3, B1 => 
                           data_in(13), B2 => n13, Y => n155);
   U85 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_14_port, A2 => n3, B1 => 
                           data_in(14), B2 => n13, Y => n153);
   U86 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_15_port, A2 => n3, B1 => 
                           data_in(15), B2 => n13, Y => n151);
   U87 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_16_port, A2 => n3, B1 => 
                           data_in(16), B2 => n11, Y => n149);
   U88 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_17_port, A2 => n3, B1 => 
                           data_in(17), B2 => n11, Y => n147);
   U89 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_18_port, A2 => n3, B1 => 
                           data_in(18), B2 => n11, Y => n145);
   U90 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_19_port, A2 => n3, B1 => 
                           data_in(19), B2 => n11, Y => n143);
   U91 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_20_port, A2 => n3, B1 => 
                           data_in(20), B2 => n11, Y => n141);
   U92 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_21_port, A2 => n3, B1 => 
                           data_in(21), B2 => n11, Y => n139);
   U93 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_22_port, A2 => n3, B1 => 
                           data_in(22), B2 => n11, Y => n137);
   U94 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_23_port, A2 => n3, B1 => 
                           data_in(23), B2 => n11, Y => n135);
   U95 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_24_port, A2 => n3, B1 => 
                           data_in(24), B2 => n11, Y => n133);
   U96 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_25_port, A2 => n3, B1 => 
                           data_in(25), B2 => n11, Y => n131);
   U97 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_26_port, A2 => n3, B1 => 
                           data_in(26), B2 => n11, Y => n129);
   U98 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_27_port, A2 => n3, B1 => 
                           data_in(27), B2 => n11, Y => n127);
   U99 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_28_port, A2 => n3, B1 => 
                           data_in(28), B2 => n9_port, Y => n125);
   U100 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_29_port, A2 => n3, B1 => 
                           data_in(29), B2 => n9_port, Y => n123);
   U101 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_30_port, A2 => n3, B1 => 
                           data_in(30), B2 => n9_port, Y => n121);
   U102 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_31_port, A2 => n3, B1 => 
                           data_in(31), B2 => n9_port, Y => n119);
   U103 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_32_port, A2 => n3, B1 => 
                           data_in(32), B2 => n9_port, Y => n117);
   U104 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_33_port, A2 => n3, B1 => 
                           data_in(33), B2 => n9_port, Y => n115);
   U105 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_34_port, A2 => n3, B1 => 
                           data_in(34), B2 => n9_port, Y => n113);
   U106 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_35_port, A2 => n3, B1 => 
                           data_in(35), B2 => n9_port, Y => n111);
   U107 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_36_port, A2 => n3, B1 => 
                           data_in(36), B2 => n9_port, Y => n109);
   U108 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_37_port, A2 => n3, B1 => 
                           data_in(37), B2 => n9_port, Y => n107);
   U109 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_38_port, A2 => n3, B1 => 
                           data_in(38), B2 => n9_port, Y => n105);
   U110 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_39_port, A2 => n3, B1 => 
                           data_in(39), B2 => n9_port, Y => n103);
   U111 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_40_port, A2 => n3, B1 => 
                           data_in(40), B2 => n7_port, Y => n101);
   U112 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_41_port, A2 => n3, B1 => 
                           data_in(41), B2 => n7_port, Y => n99);
   U113 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_42_port, A2 => n3, B1 => 
                           data_in(42), B2 => n7_port, Y => n97);
   U114 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_43_port, A2 => n3, B1 => 
                           data_in(43), B2 => n7_port, Y => n95);
   U115 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_44_port, A2 => n3, B1 => 
                           data_in(44), B2 => n7_port, Y => n93);
   U116 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_45_port, A2 => n3, B1 => 
                           data_in(45), B2 => n7_port, Y => n91);
   U117 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_46_port, A2 => n3, B1 => 
                           data_in(46), B2 => n7_port, Y => n89);
   U118 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_47_port, A2 => n3, B1 => 
                           data_in(47), B2 => n7_port, Y => n87);
   U119 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_48_port, A2 => n3, B1 => 
                           data_in(48), B2 => n7_port, Y => n85);
   U120 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_49_port, A2 => n3, B1 => 
                           data_in(49), B2 => n7_port, Y => n83);
   U121 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_50_port, A2 => n3, B1 => 
                           data_in(50), B2 => n7_port, Y => n81);
   U122 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_51_port, A2 => n3, B1 => 
                           data_in(51), B2 => n7_port, Y => n79);
   U123 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_52_port, A2 => n3, B1 => 
                           data_in(52), B2 => n5, Y => n77);
   U124 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_53_port, A2 => n3, B1 => 
                           data_in(53), B2 => n5, Y => n75);
   U125 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_54_port, A2 => n3, B1 => 
                           data_in(54), B2 => n5, Y => n73);
   U126 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_55_port, A2 => n3, B1 => 
                           data_in(55), B2 => n5, Y => n71);
   U127 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_56_port, A2 => n3, B1 => 
                           data_in(56), B2 => n5, Y => n69);
   U128 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_57_port, A2 => n3, B1 => 
                           data_in(57), B2 => n5, Y => n67);
   U129 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_58_port, A2 => n3, B1 => 
                           data_in(58), B2 => n5, Y => n65);
   U130 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_59_port, A2 => n3, B1 => 
                           data_in(59), B2 => n5, Y => n63);
   U131 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_60_port, A2 => n3, B1 => 
                           data_in(60), B2 => n5, Y => n61);
   U132 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_61_port, A2 => n3, B1 => 
                           data_in(61), B2 => n5, Y => n59);
   U133 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_62_port, A2 => n3, B1 => 
                           data_in(62), B2 => n5, Y => n57);
   U134 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_63_port, A2 => n3, B1 => 
                           data_in(63), B2 => n5, Y => n55);
   U136 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N7, Y => n236);
   U137 : OAI22xp5_ASAP7_75t_R port map( A1 => n31, A2 => read_en, B1 => n43, 
                           B2 => n45, Y => n53);
   U139 : OAI22xp5_ASAP7_75t_R port map( A1 => N9, A2 => n49, B1 => write_en, 
                           B2 => N7, Y => n51);
   write_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK 
                           => clk, RESET => n47, SET => n1, QN => N7);
   fifo_reg_1_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n55, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_63_port);
   fifo_reg_1_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n57, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_62_port);
   fifo_reg_1_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n59, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_61_port);
   fifo_reg_1_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n61, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_60_port);
   fifo_reg_0_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n171, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_63_port);
   fifo_reg_0_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n172, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_62_port);
   fifo_reg_0_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n173, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_61_port);
   fifo_reg_0_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n174, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_60_port);
   fifo_reg_1_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n167, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_3_port);
   fifo_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n168, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_2_port);
   fifo_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n169, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_1_port);
   fifo_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n170, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_0_port);
   fifo_reg_1_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n63, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_59_port);
   fifo_reg_1_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n65, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_58_port);
   fifo_reg_1_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n67, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_57_port);
   fifo_reg_1_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n69, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_56_port);
   fifo_reg_1_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n71, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_55_port);
   fifo_reg_1_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n73, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_54_port);
   fifo_reg_1_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n75, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_53_port);
   fifo_reg_1_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n77, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_52_port);
   fifo_reg_1_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_51_port);
   fifo_reg_1_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_50_port);
   fifo_reg_1_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_49_port);
   fifo_reg_1_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_48_port);
   fifo_reg_1_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_47_port);
   fifo_reg_1_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_46_port);
   fifo_reg_1_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_45_port);
   fifo_reg_1_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_44_port);
   fifo_reg_1_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_43_port);
   fifo_reg_1_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_42_port);
   fifo_reg_1_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_41_port);
   fifo_reg_1_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_40_port);
   fifo_reg_1_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_39_port);
   fifo_reg_1_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_38_port);
   fifo_reg_1_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_37_port);
   fifo_reg_1_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_36_port);
   fifo_reg_1_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_35_port);
   fifo_reg_1_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_34_port);
   fifo_reg_1_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n115, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_33_port);
   fifo_reg_1_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n117, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_32_port);
   fifo_reg_1_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n119, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_31_port);
   fifo_reg_1_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n121, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_30_port);
   fifo_reg_1_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n123, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_29_port);
   fifo_reg_1_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n125, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_28_port);
   fifo_reg_1_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n127, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_27_port);
   fifo_reg_1_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n129, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_26_port);
   fifo_reg_1_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n131, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_25_port);
   fifo_reg_1_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n133, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_24_port);
   fifo_reg_1_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n135, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_23_port);
   fifo_reg_1_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n137, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_22_port);
   fifo_reg_1_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n139, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_21_port);
   fifo_reg_1_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n141, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_20_port);
   fifo_reg_1_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n143, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_19_port);
   fifo_reg_1_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n145, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_18_port);
   fifo_reg_1_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n147, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_17_port);
   fifo_reg_1_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n149, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_16_port);
   fifo_reg_1_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n151, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_15_port);
   fifo_reg_1_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n153, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_14_port);
   fifo_reg_1_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n155, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_13_port);
   fifo_reg_1_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n157, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_12_port);
   fifo_reg_1_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n159, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_11_port);
   fifo_reg_1_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n160, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_10_port);
   fifo_reg_1_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n161, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_9_port);
   fifo_reg_1_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n162, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_8_port);
   fifo_reg_1_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n163, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_7_port);
   fifo_reg_1_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n164, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_6_port);
   fifo_reg_1_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n165, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_5_port);
   fifo_reg_1_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n166, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_4_port);
   fifo_reg_0_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n231, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_3_port);
   fifo_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n232, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_2_port);
   fifo_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n233, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_1_port);
   fifo_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n234, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_0_port);
   fifo_reg_0_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n175, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_59_port);
   fifo_reg_0_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n176, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_58_port);
   fifo_reg_0_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n177, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_57_port);
   fifo_reg_0_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n178, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_56_port);
   fifo_reg_0_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n179, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_55_port);
   fifo_reg_0_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n180, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_54_port);
   fifo_reg_0_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n181, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_53_port);
   fifo_reg_0_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n182, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_52_port);
   fifo_reg_0_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n183, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_51_port);
   fifo_reg_0_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n184, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_50_port);
   fifo_reg_0_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n185, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_49_port);
   fifo_reg_0_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n186, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_48_port);
   fifo_reg_0_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n187, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_47_port);
   fifo_reg_0_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n188, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_46_port);
   fifo_reg_0_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n189, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_45_port);
   fifo_reg_0_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n190, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_44_port);
   fifo_reg_0_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n191, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_43_port);
   fifo_reg_0_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n192, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_42_port);
   fifo_reg_0_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n193, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_41_port);
   fifo_reg_0_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n194, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_40_port);
   fifo_reg_0_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n195, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_39_port);
   fifo_reg_0_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n196, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_38_port);
   fifo_reg_0_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n197, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_37_port);
   fifo_reg_0_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n198, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_36_port);
   fifo_reg_0_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n199, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_35_port);
   fifo_reg_0_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n200, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_34_port);
   fifo_reg_0_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n201, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_33_port);
   fifo_reg_0_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n202, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_32_port);
   fifo_reg_0_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n203, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_31_port);
   fifo_reg_0_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n204, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_30_port);
   fifo_reg_0_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n205, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_29_port);
   fifo_reg_0_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n206, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_28_port);
   fifo_reg_0_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n207, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_27_port);
   fifo_reg_0_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n208, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_26_port);
   fifo_reg_0_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n209, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_25_port);
   fifo_reg_0_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n210, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_24_port);
   fifo_reg_0_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n211, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_23_port);
   fifo_reg_0_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n212, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_22_port);
   fifo_reg_0_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n213, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_21_port);
   fifo_reg_0_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n214, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_20_port);
   fifo_reg_0_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n215, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_19_port);
   fifo_reg_0_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n216, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_18_port);
   fifo_reg_0_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n217, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_17_port);
   fifo_reg_0_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n218, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_16_port);
   fifo_reg_0_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n219, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_15_port);
   fifo_reg_0_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n220, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_14_port);
   fifo_reg_0_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n221, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_13_port);
   fifo_reg_0_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n222, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_12_port);
   fifo_reg_0_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n223, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_11_port);
   fifo_reg_0_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n224, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_10_port);
   fifo_reg_0_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n225, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_9_port);
   fifo_reg_0_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n226, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_8_port);
   fifo_reg_0_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n227, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_7_port);
   fifo_reg_0_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n228, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_6_port);
   fifo_reg_0_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n229, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_5_port);
   fifo_reg_0_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n230, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_4_port);
   valid_data_reg : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n235, CLK => clk, 
                           RESET => n47, SET => n1, QN => valid_data_port);
   read_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK 
                           => clk, RESET => n47, SET => n1, QN => 
                           read_pointer_0_port);
   U69 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U135 : INVx3_ASAP7_75t_R port map( A => rst, Y => n47);
   U138 : INVx1_ASAP7_75t_R port map( A => read_en, Y => n45);
   U140 : INVx1_ASAP7_75t_R port map( A => n29, Y => n17);
   U141 : INVx1_ASAP7_75t_R port map( A => n15, Y => n3);
   U142 : INVx1_ASAP7_75t_R port map( A => n31, Y => n43);
   U207 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n29);
   U208 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n15);
   U209 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n27);
   U210 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n25);
   U211 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n23);
   U212 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n21);
   U213 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n19);
   U214 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n13);
   U215 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n11);
   U216 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n9_port);
   U217 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n7_port);
   U218 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n5);
   U219 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n31);
   U220 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n33);
   U221 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n41);
   U222 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n39);
   U223 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n37);
   U224 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n35);
   U225 : INVx1_ASAP7_75t_R port map( A => N7, Y => N9);
   U226 : INVx1_ASAP7_75t_R port map( A => write_en, Y => n49);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity fifo_buff_depth2_2 is

   port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, clk, 
         rst : in std_logic;  data_out : out std_logic_vector (63 downto 0);  
         valid_data : out std_logic);

end fifo_buff_depth2_2;

architecture SYN_rtl of fifo_buff_depth2_2 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx3_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal valid_data_port, read_pointer_0_port, fifo_1_63_port, fifo_1_62_port,
      fifo_1_61_port, fifo_1_60_port, fifo_1_59_port, fifo_1_58_port, 
      fifo_1_57_port, fifo_1_56_port, fifo_1_55_port, fifo_1_54_port, 
      fifo_1_53_port, fifo_1_52_port, fifo_1_51_port, fifo_1_50_port, 
      fifo_1_49_port, fifo_1_48_port, fifo_1_47_port, fifo_1_46_port, 
      fifo_1_45_port, fifo_1_44_port, fifo_1_43_port, fifo_1_42_port, 
      fifo_1_41_port, fifo_1_40_port, fifo_1_39_port, fifo_1_38_port, 
      fifo_1_37_port, fifo_1_36_port, fifo_1_35_port, fifo_1_34_port, 
      fifo_1_33_port, fifo_1_32_port, fifo_1_31_port, fifo_1_30_port, 
      fifo_1_29_port, fifo_1_28_port, fifo_1_27_port, fifo_1_26_port, 
      fifo_1_25_port, fifo_1_24_port, fifo_1_23_port, fifo_1_22_port, 
      fifo_1_21_port, fifo_1_20_port, fifo_1_19_port, fifo_1_18_port, 
      fifo_1_17_port, fifo_1_16_port, fifo_1_15_port, fifo_1_14_port, 
      fifo_1_13_port, fifo_1_12_port, fifo_1_11_port, fifo_1_10_port, 
      fifo_1_9_port, fifo_1_8_port, fifo_1_7_port, fifo_1_6_port, fifo_1_5_port
      , fifo_1_4_port, fifo_1_3_port, fifo_1_2_port, fifo_1_1_port, 
      fifo_1_0_port, fifo_0_63_port, fifo_0_62_port, fifo_0_61_port, 
      fifo_0_60_port, fifo_0_59_port, fifo_0_58_port, fifo_0_57_port, 
      fifo_0_56_port, fifo_0_55_port, fifo_0_54_port, fifo_0_53_port, 
      fifo_0_52_port, fifo_0_51_port, fifo_0_50_port, fifo_0_49_port, 
      fifo_0_48_port, fifo_0_47_port, fifo_0_46_port, fifo_0_45_port, 
      fifo_0_44_port, fifo_0_43_port, fifo_0_42_port, fifo_0_41_port, 
      fifo_0_40_port, fifo_0_39_port, fifo_0_38_port, fifo_0_37_port, 
      fifo_0_36_port, fifo_0_35_port, fifo_0_34_port, fifo_0_33_port, 
      fifo_0_32_port, fifo_0_31_port, fifo_0_30_port, fifo_0_29_port, 
      fifo_0_28_port, fifo_0_27_port, fifo_0_26_port, fifo_0_25_port, 
      fifo_0_24_port, fifo_0_23_port, fifo_0_22_port, fifo_0_21_port, 
      fifo_0_20_port, fifo_0_19_port, fifo_0_18_port, fifo_0_17_port, 
      fifo_0_16_port, fifo_0_15_port, fifo_0_14_port, fifo_0_13_port, 
      fifo_0_12_port, fifo_0_11_port, fifo_0_10_port, fifo_0_9_port, 
      fifo_0_8_port, fifo_0_7_port, fifo_0_6_port, fifo_0_5_port, fifo_0_4_port
      , fifo_0_3_port, fifo_0_2_port, fifo_0_1_port, fifo_0_0_port, N7, N9, n1,
      n3, n5, n7_port, n9_port, n11, n13, n15, n17, n19, n21, n23, n25, n27, 
      n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57
      , n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, 
      n87, n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, n111, 
      n113, n115, n117, n119, n121, n123, n125, n127, n129, n131, n133, n135, 
      n137, n139, n141, n143, n145, n147, n149, n151, n153, n155, n157, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238 : std_logic;

begin
   valid_data <= valid_data_port;
   
   U4 : XOR2xp5_ASAP7_75t_R port map( A => N7, B => n43, Y => n238);
   U143 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_9_port, B1 => 
                           n43, B2 => fifo_0_9_port, Y => data_out(9));
   U144 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_8_port, B1 => 
                           n43, B2 => fifo_0_8_port, Y => data_out(8));
   U145 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_7_port, B1 => 
                           n43, B2 => fifo_0_7_port, Y => data_out(7));
   U146 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_6_port, B1 => 
                           n43, B2 => fifo_0_6_port, Y => data_out(6));
   U147 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_63_port, B1 => 
                           n43, B2 => fifo_0_63_port, Y => data_out(63));
   U148 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_62_port, B1 => 
                           n43, B2 => fifo_0_62_port, Y => data_out(62));
   U149 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_61_port, B1 => 
                           n43, B2 => fifo_0_61_port, Y => data_out(61));
   U150 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_60_port, B1 => 
                           n43, B2 => fifo_0_60_port, Y => data_out(60));
   U151 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_5_port, B1 => 
                           n43, B2 => fifo_0_5_port, Y => data_out(5));
   U152 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_59_port, B1 => 
                           n43, B2 => fifo_0_59_port, Y => data_out(59));
   U153 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_58_port, B1 => 
                           n43, B2 => fifo_0_58_port, Y => data_out(58));
   U154 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_57_port, B1 => 
                           n43, B2 => fifo_0_57_port, Y => data_out(57));
   U155 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_56_port, B1 => 
                           n43, B2 => fifo_0_56_port, Y => data_out(56));
   U156 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_55_port, B1 => 
                           n43, B2 => fifo_0_55_port, Y => data_out(55));
   U157 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_54_port, B1 => 
                           n43, B2 => fifo_0_54_port, Y => data_out(54));
   U158 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_53_port, B1 => 
                           n43, B2 => fifo_0_53_port, Y => data_out(53));
   U159 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_52_port, B1 => 
                           n43, B2 => fifo_0_52_port, Y => data_out(52));
   U160 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_51_port, B1 => 
                           n43, B2 => fifo_0_51_port, Y => data_out(51));
   U161 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_50_port, B1 => 
                           n43, B2 => fifo_0_50_port, Y => data_out(50));
   U162 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_4_port, B1 => 
                           n43, B2 => fifo_0_4_port, Y => data_out(4));
   U163 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_49_port, B1 => 
                           n43, B2 => fifo_0_49_port, Y => data_out(49));
   U164 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_48_port, B1 => 
                           n43, B2 => fifo_0_48_port, Y => data_out(48));
   U165 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_47_port, B1 => 
                           n43, B2 => fifo_0_47_port, Y => data_out(47));
   U166 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_46_port, B1 => 
                           n43, B2 => fifo_0_46_port, Y => data_out(46));
   U167 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_45_port, B1 => 
                           n43, B2 => fifo_0_45_port, Y => data_out(45));
   U168 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_44_port, B1 => 
                           n43, B2 => fifo_0_44_port, Y => data_out(44));
   U169 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_43_port, B1 => 
                           n43, B2 => fifo_0_43_port, Y => data_out(43));
   U170 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_42_port, B1 => 
                           n43, B2 => fifo_0_42_port, Y => data_out(42));
   U171 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_41_port, B1 => 
                           n43, B2 => fifo_0_41_port, Y => data_out(41));
   U172 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_40_port, B1 => 
                           n43, B2 => fifo_0_40_port, Y => data_out(40));
   U173 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_3_port, B1 => 
                           n43, B2 => fifo_0_3_port, Y => data_out(3));
   U174 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_39_port, B1 => 
                           n43, B2 => fifo_0_39_port, Y => data_out(39));
   U175 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_38_port, B1 => 
                           n43, B2 => fifo_0_38_port, Y => data_out(38));
   U176 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_37_port, B1 => 
                           n43, B2 => fifo_0_37_port, Y => data_out(37));
   U177 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_36_port, B1 => 
                           n43, B2 => fifo_0_36_port, Y => data_out(36));
   U178 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_35_port, B1 => 
                           n43, B2 => fifo_0_35_port, Y => data_out(35));
   U179 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_34_port, B1 => 
                           n43, B2 => fifo_0_34_port, Y => data_out(34));
   U180 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_33_port, B1 => 
                           n43, B2 => fifo_0_33_port, Y => data_out(33));
   U181 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_32_port, B1 => 
                           n43, B2 => fifo_0_32_port, Y => data_out(32));
   U182 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_31_port, B1 => 
                           n43, B2 => fifo_0_31_port, Y => data_out(31));
   U183 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_30_port, B1 => 
                           n43, B2 => fifo_0_30_port, Y => data_out(30));
   U184 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_2_port, B1 => 
                           n43, B2 => fifo_0_2_port, Y => data_out(2));
   U185 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_29_port, B1 => 
                           n43, B2 => fifo_0_29_port, Y => data_out(29));
   U186 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_28_port, B1 => 
                           n43, B2 => fifo_0_28_port, Y => data_out(28));
   U187 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_27_port, B1 => 
                           n43, B2 => fifo_0_27_port, Y => data_out(27));
   U188 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_26_port, B1 => 
                           n43, B2 => fifo_0_26_port, Y => data_out(26));
   U189 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_25_port, B1 => 
                           n43, B2 => fifo_0_25_port, Y => data_out(25));
   U190 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_24_port, B1 => 
                           n43, B2 => fifo_0_24_port, Y => data_out(24));
   U191 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_23_port, B1 => 
                           n43, B2 => fifo_0_23_port, Y => data_out(23));
   U192 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_22_port, B1 => 
                           n43, B2 => fifo_0_22_port, Y => data_out(22));
   U193 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_21_port, B1 => 
                           n43, B2 => fifo_0_21_port, Y => data_out(21));
   U194 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_20_port, B1 => 
                           n43, B2 => fifo_0_20_port, Y => data_out(20));
   U195 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_1_port, B1 => 
                           n43, B2 => fifo_0_1_port, Y => data_out(1));
   U196 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_19_port, B1 => 
                           n43, B2 => fifo_0_19_port, Y => data_out(19));
   U197 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_18_port, B1 => 
                           n43, B2 => fifo_0_18_port, Y => data_out(18));
   U198 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_17_port, B1 => 
                           n43, B2 => fifo_0_17_port, Y => data_out(17));
   U199 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_16_port, B1 => 
                           n43, B2 => fifo_0_16_port, Y => data_out(16));
   U200 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_15_port, B1 => 
                           n43, B2 => fifo_0_15_port, Y => data_out(15));
   U201 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_14_port, B1 => 
                           n43, B2 => fifo_0_14_port, Y => data_out(14));
   U202 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_13_port, B1 => 
                           n43, B2 => fifo_0_13_port, Y => data_out(13));
   U203 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_12_port, B1 => 
                           n43, B2 => fifo_0_12_port, Y => data_out(12));
   U204 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_11_port, B1 => 
                           n43, B2 => fifo_0_11_port, Y => data_out(11));
   U205 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_10_port, B1 => 
                           n43, B2 => fifo_0_10_port, Y => data_out(10));
   U206 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_0_port, B1 => 
                           n43, B2 => fifo_0_0_port, Y => data_out(0));
   U3 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n47, A2 => n238, B => 
                           valid_data_port, C => write_en, Y => n235);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_0_port, A2 => n17, B1 => 
                           data_in(0), B2 => n29, Y => n234);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_1_port, A2 => n17, B1 => 
                           data_in(1), B2 => n29, Y => n233);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_2_port, A2 => n17, B1 => 
                           data_in(2), B2 => n29, Y => n232);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_3_port, A2 => n17, B1 => 
                           data_in(3), B2 => n29, Y => n231);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_4_port, A2 => n17, B1 => 
                           data_in(4), B2 => n27, Y => n230);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_5_port, A2 => n17, B1 => 
                           data_in(5), B2 => n27, Y => n229);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_6_port, A2 => n17, B1 => 
                           data_in(6), B2 => n27, Y => n228);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_7_port, A2 => n17, B1 => 
                           data_in(7), B2 => n27, Y => n227);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_8_port, A2 => n17, B1 => 
                           data_in(8), B2 => n27, Y => n226);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_9_port, A2 => n17, B1 => 
                           data_in(9), B2 => n27, Y => n225);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_10_port, A2 => n17, B1 => 
                           data_in(10), B2 => n27, Y => n224);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_11_port, A2 => n17, B1 => 
                           data_in(11), B2 => n27, Y => n223);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_12_port, A2 => n17, B1 => 
                           data_in(12), B2 => n27, Y => n222);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_13_port, A2 => n17, B1 => 
                           data_in(13), B2 => n27, Y => n221);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_14_port, A2 => n17, B1 => 
                           data_in(14), B2 => n27, Y => n220);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_15_port, A2 => n17, B1 => 
                           data_in(15), B2 => n27, Y => n219);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_16_port, A2 => n17, B1 => 
                           data_in(16), B2 => n25, Y => n218);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_17_port, A2 => n17, B1 => 
                           data_in(17), B2 => n25, Y => n217);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_18_port, A2 => n17, B1 => 
                           data_in(18), B2 => n25, Y => n216);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_19_port, A2 => n17, B1 => 
                           data_in(19), B2 => n25, Y => n215);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_20_port, A2 => n17, B1 => 
                           data_in(20), B2 => n25, Y => n214);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_21_port, A2 => n17, B1 => 
                           data_in(21), B2 => n25, Y => n213);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_22_port, A2 => n17, B1 => 
                           data_in(22), B2 => n25, Y => n212);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_23_port, A2 => n17, B1 => 
                           data_in(23), B2 => n25, Y => n211);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_24_port, A2 => n17, B1 => 
                           data_in(24), B2 => n25, Y => n210);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_25_port, A2 => n17, B1 => 
                           data_in(25), B2 => n25, Y => n209);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_26_port, A2 => n17, B1 => 
                           data_in(26), B2 => n25, Y => n208);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_27_port, A2 => n17, B1 => 
                           data_in(27), B2 => n25, Y => n207);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_28_port, A2 => n17, B1 => 
                           data_in(28), B2 => n23, Y => n206);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_29_port, A2 => n17, B1 => 
                           data_in(29), B2 => n23, Y => n205);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_30_port, A2 => n17, B1 => 
                           data_in(30), B2 => n23, Y => n204);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_31_port, A2 => n17, B1 => 
                           data_in(31), B2 => n23, Y => n203);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_32_port, A2 => n17, B1 => 
                           data_in(32), B2 => n23, Y => n202);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_33_port, A2 => n17, B1 => 
                           data_in(33), B2 => n23, Y => n201);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_34_port, A2 => n17, B1 => 
                           data_in(34), B2 => n23, Y => n200);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_35_port, A2 => n17, B1 => 
                           data_in(35), B2 => n23, Y => n199);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_36_port, A2 => n17, B1 => 
                           data_in(36), B2 => n23, Y => n198);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_37_port, A2 => n17, B1 => 
                           data_in(37), B2 => n23, Y => n197);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_38_port, A2 => n17, B1 => 
                           data_in(38), B2 => n23, Y => n196);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_39_port, A2 => n17, B1 => 
                           data_in(39), B2 => n23, Y => n195);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_40_port, A2 => n17, B1 => 
                           data_in(40), B2 => n21, Y => n194);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_41_port, A2 => n17, B1 => 
                           data_in(41), B2 => n21, Y => n193);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_42_port, A2 => n17, B1 => 
                           data_in(42), B2 => n21, Y => n192);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_43_port, A2 => n17, B1 => 
                           data_in(43), B2 => n21, Y => n191);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_44_port, A2 => n17, B1 => 
                           data_in(44), B2 => n21, Y => n190);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_45_port, A2 => n17, B1 => 
                           data_in(45), B2 => n21, Y => n189);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_46_port, A2 => n17, B1 => 
                           data_in(46), B2 => n21, Y => n188);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_47_port, A2 => n17, B1 => 
                           data_in(47), B2 => n21, Y => n187);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_48_port, A2 => n17, B1 => 
                           data_in(48), B2 => n21, Y => n186);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_49_port, A2 => n17, B1 => 
                           data_in(49), B2 => n21, Y => n185);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_50_port, A2 => n17, B1 => 
                           data_in(50), B2 => n21, Y => n184);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_51_port, A2 => n17, B1 => 
                           data_in(51), B2 => n21, Y => n183);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_52_port, A2 => n17, B1 => 
                           data_in(52), B2 => n19, Y => n182);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_53_port, A2 => n17, B1 => 
                           data_in(53), B2 => n19, Y => n181);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_54_port, A2 => n17, B1 => 
                           data_in(54), B2 => n19, Y => n180);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_55_port, A2 => n17, B1 => 
                           data_in(55), B2 => n19, Y => n179);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_56_port, A2 => n17, B1 => 
                           data_in(56), B2 => n19, Y => n178);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_57_port, A2 => n17, B1 => 
                           data_in(57), B2 => n19, Y => n177);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_58_port, A2 => n17, B1 => 
                           data_in(58), B2 => n19, Y => n176);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_59_port, A2 => n17, B1 => 
                           data_in(59), B2 => n19, Y => n175);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_60_port, A2 => n17, B1 => 
                           data_in(60), B2 => n19, Y => n174);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_61_port, A2 => n17, B1 => 
                           data_in(61), B2 => n19, Y => n173);
   U67 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_62_port, A2 => n17, B1 => 
                           data_in(62), B2 => n19, Y => n172);
   U68 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_63_port, A2 => n17, B1 => 
                           data_in(63), B2 => n19, Y => n171);
   U70 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N9, Y => n237);
   U71 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_0_port, A2 => n3, B1 => 
                           data_in(0), B2 => n15, Y => n170);
   U72 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_1_port, A2 => n3, B1 => 
                           data_in(1), B2 => n15, Y => n169);
   U73 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_2_port, A2 => n3, B1 => 
                           data_in(2), B2 => n15, Y => n168);
   U74 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_3_port, A2 => n3, B1 => 
                           data_in(3), B2 => n15, Y => n167);
   U75 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_4_port, A2 => n3, B1 => 
                           data_in(4), B2 => n13, Y => n166);
   U76 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_5_port, A2 => n3, B1 => 
                           data_in(5), B2 => n13, Y => n165);
   U77 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_6_port, A2 => n3, B1 => 
                           data_in(6), B2 => n13, Y => n164);
   U78 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_7_port, A2 => n3, B1 => 
                           data_in(7), B2 => n13, Y => n163);
   U79 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_8_port, A2 => n3, B1 => 
                           data_in(8), B2 => n13, Y => n162);
   U80 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_9_port, A2 => n3, B1 => 
                           data_in(9), B2 => n13, Y => n161);
   U81 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_10_port, A2 => n3, B1 => 
                           data_in(10), B2 => n13, Y => n160);
   U82 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_11_port, A2 => n3, B1 => 
                           data_in(11), B2 => n13, Y => n159);
   U83 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_12_port, A2 => n3, B1 => 
                           data_in(12), B2 => n13, Y => n157);
   U84 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_13_port, A2 => n3, B1 => 
                           data_in(13), B2 => n13, Y => n155);
   U85 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_14_port, A2 => n3, B1 => 
                           data_in(14), B2 => n13, Y => n153);
   U86 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_15_port, A2 => n3, B1 => 
                           data_in(15), B2 => n13, Y => n151);
   U87 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_16_port, A2 => n3, B1 => 
                           data_in(16), B2 => n11, Y => n149);
   U88 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_17_port, A2 => n3, B1 => 
                           data_in(17), B2 => n11, Y => n147);
   U89 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_18_port, A2 => n3, B1 => 
                           data_in(18), B2 => n11, Y => n145);
   U90 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_19_port, A2 => n3, B1 => 
                           data_in(19), B2 => n11, Y => n143);
   U91 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_20_port, A2 => n3, B1 => 
                           data_in(20), B2 => n11, Y => n141);
   U92 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_21_port, A2 => n3, B1 => 
                           data_in(21), B2 => n11, Y => n139);
   U93 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_22_port, A2 => n3, B1 => 
                           data_in(22), B2 => n11, Y => n137);
   U94 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_23_port, A2 => n3, B1 => 
                           data_in(23), B2 => n11, Y => n135);
   U95 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_24_port, A2 => n3, B1 => 
                           data_in(24), B2 => n11, Y => n133);
   U96 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_25_port, A2 => n3, B1 => 
                           data_in(25), B2 => n11, Y => n131);
   U97 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_26_port, A2 => n3, B1 => 
                           data_in(26), B2 => n11, Y => n129);
   U98 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_27_port, A2 => n3, B1 => 
                           data_in(27), B2 => n11, Y => n127);
   U99 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_28_port, A2 => n3, B1 => 
                           data_in(28), B2 => n9_port, Y => n125);
   U100 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_29_port, A2 => n3, B1 => 
                           data_in(29), B2 => n9_port, Y => n123);
   U101 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_30_port, A2 => n3, B1 => 
                           data_in(30), B2 => n9_port, Y => n121);
   U102 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_31_port, A2 => n3, B1 => 
                           data_in(31), B2 => n9_port, Y => n119);
   U103 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_32_port, A2 => n3, B1 => 
                           data_in(32), B2 => n9_port, Y => n117);
   U104 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_33_port, A2 => n3, B1 => 
                           data_in(33), B2 => n9_port, Y => n115);
   U105 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_34_port, A2 => n3, B1 => 
                           data_in(34), B2 => n9_port, Y => n113);
   U106 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_35_port, A2 => n3, B1 => 
                           data_in(35), B2 => n9_port, Y => n111);
   U107 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_36_port, A2 => n3, B1 => 
                           data_in(36), B2 => n9_port, Y => n109);
   U108 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_37_port, A2 => n3, B1 => 
                           data_in(37), B2 => n9_port, Y => n107);
   U109 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_38_port, A2 => n3, B1 => 
                           data_in(38), B2 => n9_port, Y => n105);
   U110 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_39_port, A2 => n3, B1 => 
                           data_in(39), B2 => n9_port, Y => n103);
   U111 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_40_port, A2 => n3, B1 => 
                           data_in(40), B2 => n7_port, Y => n101);
   U112 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_41_port, A2 => n3, B1 => 
                           data_in(41), B2 => n7_port, Y => n99);
   U113 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_42_port, A2 => n3, B1 => 
                           data_in(42), B2 => n7_port, Y => n97);
   U114 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_43_port, A2 => n3, B1 => 
                           data_in(43), B2 => n7_port, Y => n95);
   U115 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_44_port, A2 => n3, B1 => 
                           data_in(44), B2 => n7_port, Y => n93);
   U116 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_45_port, A2 => n3, B1 => 
                           data_in(45), B2 => n7_port, Y => n91);
   U117 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_46_port, A2 => n3, B1 => 
                           data_in(46), B2 => n7_port, Y => n89);
   U118 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_47_port, A2 => n3, B1 => 
                           data_in(47), B2 => n7_port, Y => n87);
   U119 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_48_port, A2 => n3, B1 => 
                           data_in(48), B2 => n7_port, Y => n85);
   U120 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_49_port, A2 => n3, B1 => 
                           data_in(49), B2 => n7_port, Y => n83);
   U121 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_50_port, A2 => n3, B1 => 
                           data_in(50), B2 => n7_port, Y => n81);
   U122 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_51_port, A2 => n3, B1 => 
                           data_in(51), B2 => n7_port, Y => n79);
   U123 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_52_port, A2 => n3, B1 => 
                           data_in(52), B2 => n5, Y => n77);
   U124 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_53_port, A2 => n3, B1 => 
                           data_in(53), B2 => n5, Y => n75);
   U125 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_54_port, A2 => n3, B1 => 
                           data_in(54), B2 => n5, Y => n73);
   U126 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_55_port, A2 => n3, B1 => 
                           data_in(55), B2 => n5, Y => n71);
   U127 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_56_port, A2 => n3, B1 => 
                           data_in(56), B2 => n5, Y => n69);
   U128 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_57_port, A2 => n3, B1 => 
                           data_in(57), B2 => n5, Y => n67);
   U129 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_58_port, A2 => n3, B1 => 
                           data_in(58), B2 => n5, Y => n65);
   U130 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_59_port, A2 => n3, B1 => 
                           data_in(59), B2 => n5, Y => n63);
   U131 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_60_port, A2 => n3, B1 => 
                           data_in(60), B2 => n5, Y => n61);
   U132 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_61_port, A2 => n3, B1 => 
                           data_in(61), B2 => n5, Y => n59);
   U133 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_62_port, A2 => n3, B1 => 
                           data_in(62), B2 => n5, Y => n57);
   U134 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_63_port, A2 => n3, B1 => 
                           data_in(63), B2 => n5, Y => n55);
   U136 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N7, Y => n236);
   U137 : OAI22xp5_ASAP7_75t_R port map( A1 => n31, A2 => read_en, B1 => n43, 
                           B2 => n47, Y => n53);
   U139 : OAI22xp5_ASAP7_75t_R port map( A1 => N9, A2 => n49, B1 => write_en, 
                           B2 => N7, Y => n51);
   write_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK 
                           => clk, RESET => n45, SET => n1, QN => N7);
   fifo_reg_1_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n55, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_63_port);
   fifo_reg_1_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n57, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_62_port);
   fifo_reg_1_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n59, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_61_port);
   fifo_reg_1_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n61, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_60_port);
   fifo_reg_0_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n171, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_63_port);
   fifo_reg_0_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n172, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_62_port);
   fifo_reg_0_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n173, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_61_port);
   fifo_reg_0_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n174, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_60_port);
   fifo_reg_1_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n167, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_3_port);
   fifo_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n168, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_2_port);
   fifo_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n169, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_1_port);
   fifo_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n170, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_0_port);
   fifo_reg_1_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n63, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_59_port);
   fifo_reg_1_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n65, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_58_port);
   fifo_reg_1_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n67, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_57_port);
   fifo_reg_1_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n69, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_56_port);
   fifo_reg_1_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n71, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_55_port);
   fifo_reg_1_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n73, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_54_port);
   fifo_reg_1_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n75, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_53_port);
   fifo_reg_1_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n77, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_52_port);
   fifo_reg_1_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_51_port);
   fifo_reg_1_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_50_port);
   fifo_reg_1_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_49_port);
   fifo_reg_1_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_48_port);
   fifo_reg_1_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_47_port);
   fifo_reg_1_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_46_port);
   fifo_reg_1_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_45_port);
   fifo_reg_1_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_44_port);
   fifo_reg_1_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_43_port);
   fifo_reg_1_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_42_port);
   fifo_reg_1_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_41_port);
   fifo_reg_1_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_40_port);
   fifo_reg_1_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_39_port);
   fifo_reg_1_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_38_port);
   fifo_reg_1_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_37_port);
   fifo_reg_1_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_36_port);
   fifo_reg_1_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_35_port);
   fifo_reg_1_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_34_port);
   fifo_reg_1_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n115, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_33_port);
   fifo_reg_1_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n117, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_32_port);
   fifo_reg_1_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n119, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_31_port);
   fifo_reg_1_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n121, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_30_port);
   fifo_reg_1_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n123, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_29_port);
   fifo_reg_1_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n125, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_28_port);
   fifo_reg_1_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n127, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_27_port);
   fifo_reg_1_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n129, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_26_port);
   fifo_reg_1_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n131, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_25_port);
   fifo_reg_1_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n133, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_24_port);
   fifo_reg_1_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n135, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_23_port);
   fifo_reg_1_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n137, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_22_port);
   fifo_reg_1_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n139, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_21_port);
   fifo_reg_1_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n141, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_20_port);
   fifo_reg_1_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n143, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_19_port);
   fifo_reg_1_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n145, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_18_port);
   fifo_reg_1_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n147, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_17_port);
   fifo_reg_1_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n149, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_16_port);
   fifo_reg_1_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n151, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_15_port);
   fifo_reg_1_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n153, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_14_port);
   fifo_reg_1_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n155, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_13_port);
   fifo_reg_1_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n157, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_12_port);
   fifo_reg_1_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n159, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_11_port);
   fifo_reg_1_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n160, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_10_port);
   fifo_reg_1_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n161, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_9_port);
   fifo_reg_1_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n162, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_8_port);
   fifo_reg_1_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n163, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_7_port);
   fifo_reg_1_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n164, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_6_port);
   fifo_reg_1_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n165, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_5_port);
   fifo_reg_1_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n166, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_4_port);
   fifo_reg_0_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n231, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_3_port);
   fifo_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n232, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_2_port);
   fifo_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n233, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_1_port);
   fifo_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n234, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_0_port);
   fifo_reg_0_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n175, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_59_port);
   fifo_reg_0_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n176, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_58_port);
   fifo_reg_0_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n177, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_57_port);
   fifo_reg_0_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n178, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_56_port);
   fifo_reg_0_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n179, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_55_port);
   fifo_reg_0_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n180, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_54_port);
   fifo_reg_0_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n181, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_53_port);
   fifo_reg_0_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n182, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_52_port);
   fifo_reg_0_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n183, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_51_port);
   fifo_reg_0_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n184, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_50_port);
   fifo_reg_0_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n185, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_49_port);
   fifo_reg_0_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n186, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_48_port);
   fifo_reg_0_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n187, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_47_port);
   fifo_reg_0_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n188, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_46_port);
   fifo_reg_0_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n189, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_45_port);
   fifo_reg_0_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n190, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_44_port);
   fifo_reg_0_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n191, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_43_port);
   fifo_reg_0_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n192, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_42_port);
   fifo_reg_0_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n193, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_41_port);
   fifo_reg_0_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n194, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_40_port);
   fifo_reg_0_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n195, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_39_port);
   fifo_reg_0_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n196, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_38_port);
   fifo_reg_0_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n197, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_37_port);
   fifo_reg_0_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n198, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_36_port);
   fifo_reg_0_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n199, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_35_port);
   fifo_reg_0_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n200, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_34_port);
   fifo_reg_0_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n201, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_33_port);
   fifo_reg_0_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n202, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_32_port);
   fifo_reg_0_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n203, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_31_port);
   fifo_reg_0_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n204, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_30_port);
   fifo_reg_0_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n205, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_29_port);
   fifo_reg_0_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n206, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_28_port);
   fifo_reg_0_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n207, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_27_port);
   fifo_reg_0_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n208, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_26_port);
   fifo_reg_0_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n209, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_25_port);
   fifo_reg_0_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n210, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_24_port);
   fifo_reg_0_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n211, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_23_port);
   fifo_reg_0_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n212, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_22_port);
   fifo_reg_0_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n213, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_21_port);
   fifo_reg_0_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n214, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_20_port);
   fifo_reg_0_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n215, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_19_port);
   fifo_reg_0_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n216, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_18_port);
   fifo_reg_0_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n217, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_17_port);
   fifo_reg_0_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n218, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_16_port);
   fifo_reg_0_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n219, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_15_port);
   fifo_reg_0_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n220, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_14_port);
   fifo_reg_0_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n221, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_13_port);
   fifo_reg_0_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n222, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_12_port);
   fifo_reg_0_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n223, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_11_port);
   fifo_reg_0_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n224, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_10_port);
   fifo_reg_0_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n225, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_9_port);
   fifo_reg_0_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n226, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_8_port);
   fifo_reg_0_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n227, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_7_port);
   fifo_reg_0_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n228, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_6_port);
   fifo_reg_0_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n229, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_5_port);
   fifo_reg_0_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n230, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_4_port);
   read_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK 
                           => clk, RESET => n45, SET => n1, QN => 
                           read_pointer_0_port);
   valid_data_reg : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n235, CLK => clk, 
                           RESET => n45, SET => n1, QN => valid_data_port);
   U69 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U135 : INVx3_ASAP7_75t_R port map( A => rst, Y => n45);
   U138 : INVx1_ASAP7_75t_R port map( A => n29, Y => n17);
   U140 : INVx1_ASAP7_75t_R port map( A => n15, Y => n3);
   U141 : INVx1_ASAP7_75t_R port map( A => n31, Y => n43);
   U142 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n29);
   U207 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n15);
   U208 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n27);
   U209 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n25);
   U210 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n23);
   U211 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n21);
   U212 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n19);
   U213 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n13);
   U214 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n11);
   U215 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n9_port);
   U216 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n7_port);
   U217 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n5);
   U218 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n31);
   U219 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n33);
   U220 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n41);
   U221 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n39);
   U222 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n37);
   U223 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n35);
   U224 : INVx1_ASAP7_75t_R port map( A => read_en, Y => n47);
   U225 : INVx1_ASAP7_75t_R port map( A => N7, Y => N9);
   U226 : INVx1_ASAP7_75t_R port map( A => write_en, Y => n49);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity fifo_buff_depth2_1 is

   port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, clk, 
         rst : in std_logic;  data_out : out std_logic_vector (63 downto 0);  
         valid_data : out std_logic);

end fifo_buff_depth2_1;

architecture SYN_rtl of fifo_buff_depth2_1 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx3_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal valid_data_port, read_pointer_0_port, fifo_1_63_port, fifo_1_62_port,
      fifo_1_61_port, fifo_1_60_port, fifo_1_59_port, fifo_1_58_port, 
      fifo_1_57_port, fifo_1_56_port, fifo_1_55_port, fifo_1_54_port, 
      fifo_1_53_port, fifo_1_52_port, fifo_1_51_port, fifo_1_50_port, 
      fifo_1_49_port, fifo_1_48_port, fifo_1_47_port, fifo_1_46_port, 
      fifo_1_45_port, fifo_1_44_port, fifo_1_43_port, fifo_1_42_port, 
      fifo_1_41_port, fifo_1_40_port, fifo_1_39_port, fifo_1_38_port, 
      fifo_1_37_port, fifo_1_36_port, fifo_1_35_port, fifo_1_34_port, 
      fifo_1_33_port, fifo_1_32_port, fifo_1_31_port, fifo_1_30_port, 
      fifo_1_29_port, fifo_1_28_port, fifo_1_27_port, fifo_1_26_port, 
      fifo_1_25_port, fifo_1_24_port, fifo_1_23_port, fifo_1_22_port, 
      fifo_1_21_port, fifo_1_20_port, fifo_1_19_port, fifo_1_18_port, 
      fifo_1_17_port, fifo_1_16_port, fifo_1_15_port, fifo_1_14_port, 
      fifo_1_13_port, fifo_1_12_port, fifo_1_11_port, fifo_1_10_port, 
      fifo_1_9_port, fifo_1_8_port, fifo_1_7_port, fifo_1_6_port, fifo_1_5_port
      , fifo_1_4_port, fifo_1_3_port, fifo_1_2_port, fifo_1_1_port, 
      fifo_1_0_port, fifo_0_63_port, fifo_0_62_port, fifo_0_61_port, 
      fifo_0_60_port, fifo_0_59_port, fifo_0_58_port, fifo_0_57_port, 
      fifo_0_56_port, fifo_0_55_port, fifo_0_54_port, fifo_0_53_port, 
      fifo_0_52_port, fifo_0_51_port, fifo_0_50_port, fifo_0_49_port, 
      fifo_0_48_port, fifo_0_47_port, fifo_0_46_port, fifo_0_45_port, 
      fifo_0_44_port, fifo_0_43_port, fifo_0_42_port, fifo_0_41_port, 
      fifo_0_40_port, fifo_0_39_port, fifo_0_38_port, fifo_0_37_port, 
      fifo_0_36_port, fifo_0_35_port, fifo_0_34_port, fifo_0_33_port, 
      fifo_0_32_port, fifo_0_31_port, fifo_0_30_port, fifo_0_29_port, 
      fifo_0_28_port, fifo_0_27_port, fifo_0_26_port, fifo_0_25_port, 
      fifo_0_24_port, fifo_0_23_port, fifo_0_22_port, fifo_0_21_port, 
      fifo_0_20_port, fifo_0_19_port, fifo_0_18_port, fifo_0_17_port, 
      fifo_0_16_port, fifo_0_15_port, fifo_0_14_port, fifo_0_13_port, 
      fifo_0_12_port, fifo_0_11_port, fifo_0_10_port, fifo_0_9_port, 
      fifo_0_8_port, fifo_0_7_port, fifo_0_6_port, fifo_0_5_port, fifo_0_4_port
      , fifo_0_3_port, fifo_0_2_port, fifo_0_1_port, fifo_0_0_port, N7, N9, n1,
      n3, n5, n7_port, n9_port, n11, n13, n15, n17, n19, n21, n23, n25, n27, 
      n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57
      , n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, 
      n87, n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, n111, 
      n113, n115, n117, n119, n121, n123, n125, n127, n129, n131, n133, n135, 
      n137, n139, n141, n143, n145, n147, n149, n151, n153, n155, n157, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238 : std_logic;

begin
   valid_data <= valid_data_port;
   
   U4 : XOR2xp5_ASAP7_75t_R port map( A => N7, B => n43, Y => n238);
   U143 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_9_port, B1 => 
                           n43, B2 => fifo_0_9_port, Y => data_out(9));
   U144 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_8_port, B1 => 
                           n43, B2 => fifo_0_8_port, Y => data_out(8));
   U145 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_7_port, B1 => 
                           n43, B2 => fifo_0_7_port, Y => data_out(7));
   U146 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_6_port, B1 => 
                           n43, B2 => fifo_0_6_port, Y => data_out(6));
   U147 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_63_port, B1 => 
                           n43, B2 => fifo_0_63_port, Y => data_out(63));
   U148 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_62_port, B1 => 
                           n43, B2 => fifo_0_62_port, Y => data_out(62));
   U149 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_61_port, B1 => 
                           n43, B2 => fifo_0_61_port, Y => data_out(61));
   U150 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_60_port, B1 => 
                           n43, B2 => fifo_0_60_port, Y => data_out(60));
   U151 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_5_port, B1 => 
                           n43, B2 => fifo_0_5_port, Y => data_out(5));
   U152 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_59_port, B1 => 
                           n43, B2 => fifo_0_59_port, Y => data_out(59));
   U153 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_58_port, B1 => 
                           n43, B2 => fifo_0_58_port, Y => data_out(58));
   U154 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_57_port, B1 => 
                           n43, B2 => fifo_0_57_port, Y => data_out(57));
   U155 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_56_port, B1 => 
                           n43, B2 => fifo_0_56_port, Y => data_out(56));
   U156 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_55_port, B1 => 
                           n43, B2 => fifo_0_55_port, Y => data_out(55));
   U157 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_54_port, B1 => 
                           n43, B2 => fifo_0_54_port, Y => data_out(54));
   U158 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_53_port, B1 => 
                           n43, B2 => fifo_0_53_port, Y => data_out(53));
   U159 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_52_port, B1 => 
                           n43, B2 => fifo_0_52_port, Y => data_out(52));
   U160 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_51_port, B1 => 
                           n43, B2 => fifo_0_51_port, Y => data_out(51));
   U161 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_50_port, B1 => 
                           n43, B2 => fifo_0_50_port, Y => data_out(50));
   U162 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_4_port, B1 => 
                           n43, B2 => fifo_0_4_port, Y => data_out(4));
   U163 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_49_port, B1 => 
                           n43, B2 => fifo_0_49_port, Y => data_out(49));
   U164 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_48_port, B1 => 
                           n43, B2 => fifo_0_48_port, Y => data_out(48));
   U165 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_47_port, B1 => 
                           n43, B2 => fifo_0_47_port, Y => data_out(47));
   U166 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_46_port, B1 => 
                           n43, B2 => fifo_0_46_port, Y => data_out(46));
   U167 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_45_port, B1 => 
                           n43, B2 => fifo_0_45_port, Y => data_out(45));
   U168 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_44_port, B1 => 
                           n43, B2 => fifo_0_44_port, Y => data_out(44));
   U169 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_43_port, B1 => 
                           n43, B2 => fifo_0_43_port, Y => data_out(43));
   U170 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_42_port, B1 => 
                           n43, B2 => fifo_0_42_port, Y => data_out(42));
   U171 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_41_port, B1 => 
                           n43, B2 => fifo_0_41_port, Y => data_out(41));
   U172 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_40_port, B1 => 
                           n43, B2 => fifo_0_40_port, Y => data_out(40));
   U173 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_3_port, B1 => 
                           n43, B2 => fifo_0_3_port, Y => data_out(3));
   U174 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_39_port, B1 => 
                           n43, B2 => fifo_0_39_port, Y => data_out(39));
   U175 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_38_port, B1 => 
                           n43, B2 => fifo_0_38_port, Y => data_out(38));
   U176 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_37_port, B1 => 
                           n43, B2 => fifo_0_37_port, Y => data_out(37));
   U177 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_36_port, B1 => 
                           n43, B2 => fifo_0_36_port, Y => data_out(36));
   U178 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_35_port, B1 => 
                           n43, B2 => fifo_0_35_port, Y => data_out(35));
   U179 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_34_port, B1 => 
                           n43, B2 => fifo_0_34_port, Y => data_out(34));
   U180 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_33_port, B1 => 
                           n43, B2 => fifo_0_33_port, Y => data_out(33));
   U181 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_32_port, B1 => 
                           n43, B2 => fifo_0_32_port, Y => data_out(32));
   U182 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_31_port, B1 => 
                           n43, B2 => fifo_0_31_port, Y => data_out(31));
   U183 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_30_port, B1 => 
                           n43, B2 => fifo_0_30_port, Y => data_out(30));
   U184 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_2_port, B1 => 
                           n43, B2 => fifo_0_2_port, Y => data_out(2));
   U185 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_29_port, B1 => 
                           n43, B2 => fifo_0_29_port, Y => data_out(29));
   U186 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_28_port, B1 => 
                           n43, B2 => fifo_0_28_port, Y => data_out(28));
   U187 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_27_port, B1 => 
                           n43, B2 => fifo_0_27_port, Y => data_out(27));
   U188 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_26_port, B1 => 
                           n43, B2 => fifo_0_26_port, Y => data_out(26));
   U189 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_25_port, B1 => 
                           n43, B2 => fifo_0_25_port, Y => data_out(25));
   U190 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_24_port, B1 => 
                           n43, B2 => fifo_0_24_port, Y => data_out(24));
   U191 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_23_port, B1 => 
                           n43, B2 => fifo_0_23_port, Y => data_out(23));
   U192 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_22_port, B1 => 
                           n43, B2 => fifo_0_22_port, Y => data_out(22));
   U193 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_21_port, B1 => 
                           n43, B2 => fifo_0_21_port, Y => data_out(21));
   U194 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_20_port, B1 => 
                           n43, B2 => fifo_0_20_port, Y => data_out(20));
   U195 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_1_port, B1 => 
                           n43, B2 => fifo_0_1_port, Y => data_out(1));
   U196 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_19_port, B1 => 
                           n43, B2 => fifo_0_19_port, Y => data_out(19));
   U197 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_18_port, B1 => 
                           n43, B2 => fifo_0_18_port, Y => data_out(18));
   U198 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_17_port, B1 => 
                           n43, B2 => fifo_0_17_port, Y => data_out(17));
   U199 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_16_port, B1 => 
                           n43, B2 => fifo_0_16_port, Y => data_out(16));
   U200 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_15_port, B1 => 
                           n43, B2 => fifo_0_15_port, Y => data_out(15));
   U201 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_14_port, B1 => 
                           n43, B2 => fifo_0_14_port, Y => data_out(14));
   U202 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_13_port, B1 => 
                           n43, B2 => fifo_0_13_port, Y => data_out(13));
   U203 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_12_port, B1 => 
                           n43, B2 => fifo_0_12_port, Y => data_out(12));
   U204 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_11_port, B1 => 
                           n43, B2 => fifo_0_11_port, Y => data_out(11));
   U205 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_10_port, B1 => 
                           n43, B2 => fifo_0_10_port, Y => data_out(10));
   U206 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_0_port, B1 => 
                           n43, B2 => fifo_0_0_port, Y => data_out(0));
   U3 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n45, A2 => n238, B => 
                           valid_data_port, C => write_en, Y => n235);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_0_port, A2 => n17, B1 => 
                           data_in(0), B2 => n29, Y => n234);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_1_port, A2 => n17, B1 => 
                           data_in(1), B2 => n29, Y => n233);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_2_port, A2 => n17, B1 => 
                           data_in(2), B2 => n29, Y => n232);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_3_port, A2 => n17, B1 => 
                           data_in(3), B2 => n29, Y => n231);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_4_port, A2 => n17, B1 => 
                           data_in(4), B2 => n27, Y => n230);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_5_port, A2 => n17, B1 => 
                           data_in(5), B2 => n27, Y => n229);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_6_port, A2 => n17, B1 => 
                           data_in(6), B2 => n27, Y => n228);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_7_port, A2 => n17, B1 => 
                           data_in(7), B2 => n27, Y => n227);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_8_port, A2 => n17, B1 => 
                           data_in(8), B2 => n27, Y => n226);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_9_port, A2 => n17, B1 => 
                           data_in(9), B2 => n27, Y => n225);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_10_port, A2 => n17, B1 => 
                           data_in(10), B2 => n27, Y => n224);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_11_port, A2 => n17, B1 => 
                           data_in(11), B2 => n27, Y => n223);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_12_port, A2 => n17, B1 => 
                           data_in(12), B2 => n27, Y => n222);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_13_port, A2 => n17, B1 => 
                           data_in(13), B2 => n27, Y => n221);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_14_port, A2 => n17, B1 => 
                           data_in(14), B2 => n27, Y => n220);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_15_port, A2 => n17, B1 => 
                           data_in(15), B2 => n27, Y => n219);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_16_port, A2 => n17, B1 => 
                           data_in(16), B2 => n25, Y => n218);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_17_port, A2 => n17, B1 => 
                           data_in(17), B2 => n25, Y => n217);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_18_port, A2 => n17, B1 => 
                           data_in(18), B2 => n25, Y => n216);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_19_port, A2 => n17, B1 => 
                           data_in(19), B2 => n25, Y => n215);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_20_port, A2 => n17, B1 => 
                           data_in(20), B2 => n25, Y => n214);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_21_port, A2 => n17, B1 => 
                           data_in(21), B2 => n25, Y => n213);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_22_port, A2 => n17, B1 => 
                           data_in(22), B2 => n25, Y => n212);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_23_port, A2 => n17, B1 => 
                           data_in(23), B2 => n25, Y => n211);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_24_port, A2 => n17, B1 => 
                           data_in(24), B2 => n25, Y => n210);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_25_port, A2 => n17, B1 => 
                           data_in(25), B2 => n25, Y => n209);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_26_port, A2 => n17, B1 => 
                           data_in(26), B2 => n25, Y => n208);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_27_port, A2 => n17, B1 => 
                           data_in(27), B2 => n25, Y => n207);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_28_port, A2 => n17, B1 => 
                           data_in(28), B2 => n23, Y => n206);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_29_port, A2 => n17, B1 => 
                           data_in(29), B2 => n23, Y => n205);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_30_port, A2 => n17, B1 => 
                           data_in(30), B2 => n23, Y => n204);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_31_port, A2 => n17, B1 => 
                           data_in(31), B2 => n23, Y => n203);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_32_port, A2 => n17, B1 => 
                           data_in(32), B2 => n23, Y => n202);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_33_port, A2 => n17, B1 => 
                           data_in(33), B2 => n23, Y => n201);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_34_port, A2 => n17, B1 => 
                           data_in(34), B2 => n23, Y => n200);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_35_port, A2 => n17, B1 => 
                           data_in(35), B2 => n23, Y => n199);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_36_port, A2 => n17, B1 => 
                           data_in(36), B2 => n23, Y => n198);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_37_port, A2 => n17, B1 => 
                           data_in(37), B2 => n23, Y => n197);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_38_port, A2 => n17, B1 => 
                           data_in(38), B2 => n23, Y => n196);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_39_port, A2 => n17, B1 => 
                           data_in(39), B2 => n23, Y => n195);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_40_port, A2 => n17, B1 => 
                           data_in(40), B2 => n21, Y => n194);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_41_port, A2 => n17, B1 => 
                           data_in(41), B2 => n21, Y => n193);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_42_port, A2 => n17, B1 => 
                           data_in(42), B2 => n21, Y => n192);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_43_port, A2 => n17, B1 => 
                           data_in(43), B2 => n21, Y => n191);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_44_port, A2 => n17, B1 => 
                           data_in(44), B2 => n21, Y => n190);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_45_port, A2 => n17, B1 => 
                           data_in(45), B2 => n21, Y => n189);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_46_port, A2 => n17, B1 => 
                           data_in(46), B2 => n21, Y => n188);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_47_port, A2 => n17, B1 => 
                           data_in(47), B2 => n21, Y => n187);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_48_port, A2 => n17, B1 => 
                           data_in(48), B2 => n21, Y => n186);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_49_port, A2 => n17, B1 => 
                           data_in(49), B2 => n21, Y => n185);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_50_port, A2 => n17, B1 => 
                           data_in(50), B2 => n21, Y => n184);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_51_port, A2 => n17, B1 => 
                           data_in(51), B2 => n21, Y => n183);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_52_port, A2 => n17, B1 => 
                           data_in(52), B2 => n19, Y => n182);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_53_port, A2 => n17, B1 => 
                           data_in(53), B2 => n19, Y => n181);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_54_port, A2 => n17, B1 => 
                           data_in(54), B2 => n19, Y => n180);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_55_port, A2 => n17, B1 => 
                           data_in(55), B2 => n19, Y => n179);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_56_port, A2 => n17, B1 => 
                           data_in(56), B2 => n19, Y => n178);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_57_port, A2 => n17, B1 => 
                           data_in(57), B2 => n19, Y => n177);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_58_port, A2 => n17, B1 => 
                           data_in(58), B2 => n19, Y => n176);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_59_port, A2 => n17, B1 => 
                           data_in(59), B2 => n19, Y => n175);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_60_port, A2 => n17, B1 => 
                           data_in(60), B2 => n19, Y => n174);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_61_port, A2 => n17, B1 => 
                           data_in(61), B2 => n19, Y => n173);
   U67 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_62_port, A2 => n17, B1 => 
                           data_in(62), B2 => n19, Y => n172);
   U68 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_63_port, A2 => n17, B1 => 
                           data_in(63), B2 => n19, Y => n171);
   U70 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N9, Y => n237);
   U71 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_0_port, A2 => n3, B1 => 
                           data_in(0), B2 => n15, Y => n170);
   U72 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_1_port, A2 => n3, B1 => 
                           data_in(1), B2 => n15, Y => n169);
   U73 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_2_port, A2 => n3, B1 => 
                           data_in(2), B2 => n15, Y => n168);
   U74 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_3_port, A2 => n3, B1 => 
                           data_in(3), B2 => n15, Y => n167);
   U75 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_4_port, A2 => n3, B1 => 
                           data_in(4), B2 => n13, Y => n166);
   U76 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_5_port, A2 => n3, B1 => 
                           data_in(5), B2 => n13, Y => n165);
   U77 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_6_port, A2 => n3, B1 => 
                           data_in(6), B2 => n13, Y => n164);
   U78 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_7_port, A2 => n3, B1 => 
                           data_in(7), B2 => n13, Y => n163);
   U79 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_8_port, A2 => n3, B1 => 
                           data_in(8), B2 => n13, Y => n162);
   U80 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_9_port, A2 => n3, B1 => 
                           data_in(9), B2 => n13, Y => n161);
   U81 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_10_port, A2 => n3, B1 => 
                           data_in(10), B2 => n13, Y => n160);
   U82 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_11_port, A2 => n3, B1 => 
                           data_in(11), B2 => n13, Y => n159);
   U83 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_12_port, A2 => n3, B1 => 
                           data_in(12), B2 => n13, Y => n157);
   U84 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_13_port, A2 => n3, B1 => 
                           data_in(13), B2 => n13, Y => n155);
   U85 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_14_port, A2 => n3, B1 => 
                           data_in(14), B2 => n13, Y => n153);
   U86 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_15_port, A2 => n3, B1 => 
                           data_in(15), B2 => n13, Y => n151);
   U87 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_16_port, A2 => n3, B1 => 
                           data_in(16), B2 => n11, Y => n149);
   U88 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_17_port, A2 => n3, B1 => 
                           data_in(17), B2 => n11, Y => n147);
   U89 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_18_port, A2 => n3, B1 => 
                           data_in(18), B2 => n11, Y => n145);
   U90 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_19_port, A2 => n3, B1 => 
                           data_in(19), B2 => n11, Y => n143);
   U91 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_20_port, A2 => n3, B1 => 
                           data_in(20), B2 => n11, Y => n141);
   U92 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_21_port, A2 => n3, B1 => 
                           data_in(21), B2 => n11, Y => n139);
   U93 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_22_port, A2 => n3, B1 => 
                           data_in(22), B2 => n11, Y => n137);
   U94 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_23_port, A2 => n3, B1 => 
                           data_in(23), B2 => n11, Y => n135);
   U95 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_24_port, A2 => n3, B1 => 
                           data_in(24), B2 => n11, Y => n133);
   U96 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_25_port, A2 => n3, B1 => 
                           data_in(25), B2 => n11, Y => n131);
   U97 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_26_port, A2 => n3, B1 => 
                           data_in(26), B2 => n11, Y => n129);
   U98 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_27_port, A2 => n3, B1 => 
                           data_in(27), B2 => n11, Y => n127);
   U99 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_28_port, A2 => n3, B1 => 
                           data_in(28), B2 => n9_port, Y => n125);
   U100 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_29_port, A2 => n3, B1 => 
                           data_in(29), B2 => n9_port, Y => n123);
   U101 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_30_port, A2 => n3, B1 => 
                           data_in(30), B2 => n9_port, Y => n121);
   U102 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_31_port, A2 => n3, B1 => 
                           data_in(31), B2 => n9_port, Y => n119);
   U103 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_32_port, A2 => n3, B1 => 
                           data_in(32), B2 => n9_port, Y => n117);
   U104 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_33_port, A2 => n3, B1 => 
                           data_in(33), B2 => n9_port, Y => n115);
   U105 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_34_port, A2 => n3, B1 => 
                           data_in(34), B2 => n9_port, Y => n113);
   U106 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_35_port, A2 => n3, B1 => 
                           data_in(35), B2 => n9_port, Y => n111);
   U107 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_36_port, A2 => n3, B1 => 
                           data_in(36), B2 => n9_port, Y => n109);
   U108 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_37_port, A2 => n3, B1 => 
                           data_in(37), B2 => n9_port, Y => n107);
   U109 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_38_port, A2 => n3, B1 => 
                           data_in(38), B2 => n9_port, Y => n105);
   U110 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_39_port, A2 => n3, B1 => 
                           data_in(39), B2 => n9_port, Y => n103);
   U111 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_40_port, A2 => n3, B1 => 
                           data_in(40), B2 => n7_port, Y => n101);
   U112 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_41_port, A2 => n3, B1 => 
                           data_in(41), B2 => n7_port, Y => n99);
   U113 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_42_port, A2 => n3, B1 => 
                           data_in(42), B2 => n7_port, Y => n97);
   U114 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_43_port, A2 => n3, B1 => 
                           data_in(43), B2 => n7_port, Y => n95);
   U115 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_44_port, A2 => n3, B1 => 
                           data_in(44), B2 => n7_port, Y => n93);
   U116 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_45_port, A2 => n3, B1 => 
                           data_in(45), B2 => n7_port, Y => n91);
   U117 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_46_port, A2 => n3, B1 => 
                           data_in(46), B2 => n7_port, Y => n89);
   U118 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_47_port, A2 => n3, B1 => 
                           data_in(47), B2 => n7_port, Y => n87);
   U119 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_48_port, A2 => n3, B1 => 
                           data_in(48), B2 => n7_port, Y => n85);
   U120 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_49_port, A2 => n3, B1 => 
                           data_in(49), B2 => n7_port, Y => n83);
   U121 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_50_port, A2 => n3, B1 => 
                           data_in(50), B2 => n7_port, Y => n81);
   U122 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_51_port, A2 => n3, B1 => 
                           data_in(51), B2 => n7_port, Y => n79);
   U123 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_52_port, A2 => n3, B1 => 
                           data_in(52), B2 => n5, Y => n77);
   U124 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_53_port, A2 => n3, B1 => 
                           data_in(53), B2 => n5, Y => n75);
   U125 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_54_port, A2 => n3, B1 => 
                           data_in(54), B2 => n5, Y => n73);
   U126 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_55_port, A2 => n3, B1 => 
                           data_in(55), B2 => n5, Y => n71);
   U127 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_56_port, A2 => n3, B1 => 
                           data_in(56), B2 => n5, Y => n69);
   U128 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_57_port, A2 => n3, B1 => 
                           data_in(57), B2 => n5, Y => n67);
   U129 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_58_port, A2 => n3, B1 => 
                           data_in(58), B2 => n5, Y => n65);
   U130 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_59_port, A2 => n3, B1 => 
                           data_in(59), B2 => n5, Y => n63);
   U131 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_60_port, A2 => n3, B1 => 
                           data_in(60), B2 => n5, Y => n61);
   U132 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_61_port, A2 => n3, B1 => 
                           data_in(61), B2 => n5, Y => n59);
   U133 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_62_port, A2 => n3, B1 => 
                           data_in(62), B2 => n5, Y => n57);
   U134 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_63_port, A2 => n3, B1 => 
                           data_in(63), B2 => n5, Y => n55);
   U136 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N7, Y => n236);
   U137 : OAI22xp5_ASAP7_75t_R port map( A1 => n31, A2 => read_en, B1 => n43, 
                           B2 => n45, Y => n53);
   U139 : OAI22xp5_ASAP7_75t_R port map( A1 => N9, A2 => n49, B1 => write_en, 
                           B2 => N7, Y => n51);
   write_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK 
                           => clk, RESET => n47, SET => n1, QN => N7);
   fifo_reg_1_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n55, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_63_port);
   fifo_reg_1_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n57, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_62_port);
   fifo_reg_1_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n59, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_61_port);
   fifo_reg_1_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n61, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_60_port);
   fifo_reg_0_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n171, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_63_port);
   fifo_reg_0_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n172, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_62_port);
   fifo_reg_0_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n173, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_61_port);
   fifo_reg_0_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n174, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_60_port);
   fifo_reg_1_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n167, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_3_port);
   fifo_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n168, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_2_port);
   fifo_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n169, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_1_port);
   fifo_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n170, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_0_port);
   fifo_reg_1_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n63, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_59_port);
   fifo_reg_1_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n65, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_58_port);
   fifo_reg_1_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n67, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_57_port);
   fifo_reg_1_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n69, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_56_port);
   fifo_reg_1_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n71, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_55_port);
   fifo_reg_1_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n73, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_54_port);
   fifo_reg_1_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n75, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_53_port);
   fifo_reg_1_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n77, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_52_port);
   fifo_reg_1_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_51_port);
   fifo_reg_1_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_50_port);
   fifo_reg_1_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_49_port);
   fifo_reg_1_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_48_port);
   fifo_reg_1_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_47_port);
   fifo_reg_1_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_46_port);
   fifo_reg_1_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_45_port);
   fifo_reg_1_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_44_port);
   fifo_reg_1_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_43_port);
   fifo_reg_1_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_42_port);
   fifo_reg_1_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_41_port);
   fifo_reg_1_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_40_port);
   fifo_reg_1_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_39_port);
   fifo_reg_1_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_38_port);
   fifo_reg_1_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_37_port);
   fifo_reg_1_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_36_port);
   fifo_reg_1_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_35_port);
   fifo_reg_1_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_34_port);
   fifo_reg_1_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n115, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_33_port);
   fifo_reg_1_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n117, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_32_port);
   fifo_reg_1_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n119, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_31_port);
   fifo_reg_1_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n121, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_30_port);
   fifo_reg_1_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n123, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_29_port);
   fifo_reg_1_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n125, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_28_port);
   fifo_reg_1_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n127, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_27_port);
   fifo_reg_1_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n129, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_26_port);
   fifo_reg_1_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n131, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_25_port);
   fifo_reg_1_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n133, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_24_port);
   fifo_reg_1_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n135, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_23_port);
   fifo_reg_1_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n137, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_22_port);
   fifo_reg_1_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n139, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_21_port);
   fifo_reg_1_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n141, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_20_port);
   fifo_reg_1_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n143, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_19_port);
   fifo_reg_1_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n145, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_18_port);
   fifo_reg_1_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n147, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_17_port);
   fifo_reg_1_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n149, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_16_port);
   fifo_reg_1_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n151, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_15_port);
   fifo_reg_1_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n153, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_14_port);
   fifo_reg_1_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n155, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_13_port);
   fifo_reg_1_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n157, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_12_port);
   fifo_reg_1_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n159, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_11_port);
   fifo_reg_1_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n160, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_1_10_port);
   fifo_reg_1_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n161, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_9_port);
   fifo_reg_1_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n162, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_8_port);
   fifo_reg_1_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n163, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_7_port);
   fifo_reg_1_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n164, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_6_port);
   fifo_reg_1_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n165, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_5_port);
   fifo_reg_1_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n166, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_1_4_port);
   fifo_reg_0_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n231, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_3_port);
   fifo_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n232, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_2_port);
   fifo_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n233, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_1_port);
   fifo_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n234, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_0_port);
   fifo_reg_0_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n175, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_59_port);
   fifo_reg_0_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n176, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_58_port);
   fifo_reg_0_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n177, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_57_port);
   fifo_reg_0_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n178, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_56_port);
   fifo_reg_0_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n179, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_55_port);
   fifo_reg_0_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n180, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_54_port);
   fifo_reg_0_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n181, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_53_port);
   fifo_reg_0_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n182, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_52_port);
   fifo_reg_0_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n183, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_51_port);
   fifo_reg_0_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n184, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_50_port);
   fifo_reg_0_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n185, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_49_port);
   fifo_reg_0_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n186, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_48_port);
   fifo_reg_0_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n187, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_47_port);
   fifo_reg_0_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n188, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_46_port);
   fifo_reg_0_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n189, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_45_port);
   fifo_reg_0_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n190, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_44_port);
   fifo_reg_0_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n191, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_43_port);
   fifo_reg_0_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n192, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_42_port);
   fifo_reg_0_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n193, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_41_port);
   fifo_reg_0_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n194, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_40_port);
   fifo_reg_0_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n195, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_39_port);
   fifo_reg_0_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n196, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_38_port);
   fifo_reg_0_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n197, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_37_port);
   fifo_reg_0_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n198, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_36_port);
   fifo_reg_0_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n199, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_35_port);
   fifo_reg_0_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n200, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_34_port);
   fifo_reg_0_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n201, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_33_port);
   fifo_reg_0_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n202, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_32_port);
   fifo_reg_0_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n203, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_31_port);
   fifo_reg_0_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n204, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_30_port);
   fifo_reg_0_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n205, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_29_port);
   fifo_reg_0_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n206, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_28_port);
   fifo_reg_0_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n207, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_27_port);
   fifo_reg_0_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n208, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_26_port);
   fifo_reg_0_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n209, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_25_port);
   fifo_reg_0_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n210, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_24_port);
   fifo_reg_0_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n211, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_23_port);
   fifo_reg_0_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n212, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_22_port);
   fifo_reg_0_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n213, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_21_port);
   fifo_reg_0_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n214, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_20_port);
   fifo_reg_0_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n215, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_19_port);
   fifo_reg_0_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n216, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_18_port);
   fifo_reg_0_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n217, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_17_port);
   fifo_reg_0_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n218, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_16_port);
   fifo_reg_0_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n219, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_15_port);
   fifo_reg_0_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n220, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_14_port);
   fifo_reg_0_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n221, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_13_port);
   fifo_reg_0_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n222, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_12_port);
   fifo_reg_0_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n223, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_11_port);
   fifo_reg_0_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n224, CLK => 
                           clk, RESET => n47, SET => n1, QN => fifo_0_10_port);
   fifo_reg_0_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n225, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_9_port);
   fifo_reg_0_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n226, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_8_port);
   fifo_reg_0_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n227, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_7_port);
   fifo_reg_0_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n228, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_6_port);
   fifo_reg_0_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n229, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_5_port);
   fifo_reg_0_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n230, CLK => clk
                           , RESET => n47, SET => n1, QN => fifo_0_4_port);
   valid_data_reg : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n235, CLK => clk, 
                           RESET => n47, SET => n1, QN => valid_data_port);
   read_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK 
                           => clk, RESET => n47, SET => n1, QN => 
                           read_pointer_0_port);
   U69 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U135 : INVx3_ASAP7_75t_R port map( A => rst, Y => n47);
   U138 : INVx1_ASAP7_75t_R port map( A => read_en, Y => n45);
   U140 : INVx1_ASAP7_75t_R port map( A => n29, Y => n17);
   U141 : INVx1_ASAP7_75t_R port map( A => n15, Y => n3);
   U142 : INVx1_ASAP7_75t_R port map( A => n31, Y => n43);
   U207 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n29);
   U208 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n15);
   U209 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n27);
   U210 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n25);
   U211 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n23);
   U212 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n21);
   U213 : HB1xp67_ASAP7_75t_R port map( A => n237, Y => n19);
   U214 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n13);
   U215 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n11);
   U216 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n9_port);
   U217 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n7_port);
   U218 : HB1xp67_ASAP7_75t_R port map( A => n236, Y => n5);
   U219 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n31);
   U220 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n33);
   U221 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n41);
   U222 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n39);
   U223 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n37);
   U224 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n35);
   U225 : INVx1_ASAP7_75t_R port map( A => N7, Y => N9);
   U226 : INVx1_ASAP7_75t_R port map( A => write_en, Y => n49);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity output_register_vc_num2_vc_num_out2_5 is

   port( clk, rst : in std_logic;  data_tx : in std_logic_vector (63 downto 0);
         vc_write_tx, incr_tx : in std_logic_vector (1 downto 0);  data_tx_pl :
         out std_logic_vector (63 downto 0);  vc_write_tx_pl, incr_tx_pl : out 
         std_logic_vector (1 downto 0));

end output_register_vc_num2_vc_num_out2_5;

architecture SYN_rtl of output_register_vc_num2_vc_num_out2_5 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx2_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal data_tx_pl_63_port, data_tx_pl_62_port, data_tx_pl_61_port, 
      data_tx_pl_60_port, data_tx_pl_59_port, data_tx_pl_58_port, 
      data_tx_pl_57_port, data_tx_pl_56_port, data_tx_pl_55_port, 
      data_tx_pl_54_port, data_tx_pl_53_port, data_tx_pl_52_port, 
      data_tx_pl_51_port, data_tx_pl_50_port, data_tx_pl_49_port, 
      data_tx_pl_48_port, data_tx_pl_47_port, data_tx_pl_46_port, 
      data_tx_pl_45_port, data_tx_pl_44_port, data_tx_pl_43_port, 
      data_tx_pl_42_port, data_tx_pl_41_port, data_tx_pl_40_port, 
      data_tx_pl_39_port, data_tx_pl_38_port, data_tx_pl_37_port, 
      data_tx_pl_36_port, data_tx_pl_35_port, data_tx_pl_34_port, 
      data_tx_pl_33_port, data_tx_pl_32_port, data_tx_pl_31_port, 
      data_tx_pl_30_port, data_tx_pl_29_port, data_tx_pl_28_port, 
      data_tx_pl_27_port, data_tx_pl_26_port, data_tx_pl_25_port, 
      data_tx_pl_24_port, data_tx_pl_23_port, data_tx_pl_22_port, 
      data_tx_pl_21_port, data_tx_pl_20_port, data_tx_pl_19_port, 
      data_tx_pl_18_port, data_tx_pl_17_port, data_tx_pl_16_port, 
      data_tx_pl_15_port, data_tx_pl_14_port, data_tx_pl_13_port, 
      data_tx_pl_12_port, data_tx_pl_11_port, data_tx_pl_10_port, 
      data_tx_pl_9_port, data_tx_pl_8_port, data_tx_pl_7_port, 
      data_tx_pl_6_port, data_tx_pl_5_port, data_tx_pl_4_port, 
      data_tx_pl_3_port, data_tx_pl_2_port, data_tx_pl_1_port, 
      data_tx_pl_0_port, n1, n3, n4, n5, n6, n8, n10, n12, n14, n16, n18, n20, 
      n22, n24, n26, n28, n30, n32, n34, n36, n38, n40, n42, n44, n46, n48, n50
      , n52, n54, n56, n58, n60, n62, n64, n66, n68, n70, n72, n74, n76, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
      n107, n108, n109, n110, n111, n112, n113, n114, n115 : std_logic;

begin
   data_tx_pl <= ( data_tx_pl_63_port, data_tx_pl_62_port, data_tx_pl_61_port, 
      data_tx_pl_60_port, data_tx_pl_59_port, data_tx_pl_58_port, 
      data_tx_pl_57_port, data_tx_pl_56_port, data_tx_pl_55_port, 
      data_tx_pl_54_port, data_tx_pl_53_port, data_tx_pl_52_port, 
      data_tx_pl_51_port, data_tx_pl_50_port, data_tx_pl_49_port, 
      data_tx_pl_48_port, data_tx_pl_47_port, data_tx_pl_46_port, 
      data_tx_pl_45_port, data_tx_pl_44_port, data_tx_pl_43_port, 
      data_tx_pl_42_port, data_tx_pl_41_port, data_tx_pl_40_port, 
      data_tx_pl_39_port, data_tx_pl_38_port, data_tx_pl_37_port, 
      data_tx_pl_36_port, data_tx_pl_35_port, data_tx_pl_34_port, 
      data_tx_pl_33_port, data_tx_pl_32_port, data_tx_pl_31_port, 
      data_tx_pl_30_port, data_tx_pl_29_port, data_tx_pl_28_port, 
      data_tx_pl_27_port, data_tx_pl_26_port, data_tx_pl_25_port, 
      data_tx_pl_24_port, data_tx_pl_23_port, data_tx_pl_22_port, 
      data_tx_pl_21_port, data_tx_pl_20_port, data_tx_pl_19_port, 
      data_tx_pl_18_port, data_tx_pl_17_port, data_tx_pl_16_port, 
      data_tx_pl_15_port, data_tx_pl_14_port, data_tx_pl_13_port, 
      data_tx_pl_12_port, data_tx_pl_11_port, data_tx_pl_10_port, 
      data_tx_pl_9_port, data_tx_pl_8_port, data_tx_pl_7_port, 
      data_tx_pl_6_port, data_tx_pl_5_port, data_tx_pl_4_port, 
      data_tx_pl_3_port, data_tx_pl_2_port, data_tx_pl_1_port, 
      data_tx_pl_0_port );
   
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(0), A2 => n3, B1 => 
                           data_tx_pl_0_port, B2 => n12, Y => n114);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(1), A2 => n3, B1 => 
                           data_tx_pl_1_port, B2 => n12, Y => n113);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(2), A2 => n3, B1 => 
                           data_tx_pl_2_port, B2 => n12, Y => n112);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(3), A2 => n3, B1 => 
                           data_tx_pl_3_port, B2 => n12, Y => n111);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(4), A2 => n3, B1 => 
                           data_tx_pl_4_port, B2 => n10, Y => n110);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(5), A2 => n3, B1 => 
                           data_tx_pl_5_port, B2 => n10, Y => n109);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(6), A2 => n3, B1 => 
                           data_tx_pl_6_port, B2 => n10, Y => n108);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(7), A2 => n3, B1 => 
                           data_tx_pl_7_port, B2 => n10, Y => n107);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(8), A2 => n3, B1 => 
                           data_tx_pl_8_port, B2 => n10, Y => n106);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(9), A2 => n3, B1 => 
                           data_tx_pl_9_port, B2 => n10, Y => n105);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(10), A2 => n3, B1 => 
                           data_tx_pl_10_port, B2 => n10, Y => n104);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(11), A2 => n3, B1 => 
                           data_tx_pl_11_port, B2 => n10, Y => n103);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(12), A2 => n3, B1 => 
                           data_tx_pl_12_port, B2 => n10, Y => n102);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(13), A2 => n3, B1 => 
                           data_tx_pl_13_port, B2 => n10, Y => n101);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(14), A2 => n3, B1 => 
                           data_tx_pl_14_port, B2 => n10, Y => n100);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(15), A2 => n3, B1 => 
                           data_tx_pl_15_port, B2 => n10, Y => n99);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(16), A2 => n3, B1 => 
                           data_tx_pl_16_port, B2 => n8, Y => n98);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(17), A2 => n3, B1 => 
                           data_tx_pl_17_port, B2 => n8, Y => n97);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(18), A2 => n3, B1 => 
                           data_tx_pl_18_port, B2 => n8, Y => n96);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(19), A2 => n3, B1 => 
                           data_tx_pl_19_port, B2 => n8, Y => n95);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(20), A2 => n3, B1 => 
                           data_tx_pl_20_port, B2 => n8, Y => n94);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(21), A2 => n3, B1 => 
                           data_tx_pl_21_port, B2 => n8, Y => n93);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(22), A2 => n3, B1 => 
                           data_tx_pl_22_port, B2 => n8, Y => n92);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(23), A2 => n3, B1 => 
                           data_tx_pl_23_port, B2 => n8, Y => n91);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(24), A2 => n3, B1 => 
                           data_tx_pl_24_port, B2 => n8, Y => n90);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(25), A2 => n3, B1 => 
                           data_tx_pl_25_port, B2 => n8, Y => n89);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(26), A2 => n3, B1 => 
                           data_tx_pl_26_port, B2 => n8, Y => n88);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(27), A2 => n3, B1 => 
                           data_tx_pl_27_port, B2 => n8, Y => n87);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(28), A2 => n3, B1 => 
                           data_tx_pl_28_port, B2 => n6, Y => n86);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(29), A2 => n3, B1 => 
                           data_tx_pl_29_port, B2 => n6, Y => n85);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(30), A2 => n3, B1 => 
                           data_tx_pl_30_port, B2 => n6, Y => n84);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(31), A2 => n3, B1 => 
                           data_tx_pl_31_port, B2 => n6, Y => n83);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(32), A2 => n3, B1 => 
                           data_tx_pl_32_port, B2 => n6, Y => n82);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(33), A2 => n3, B1 => 
                           data_tx_pl_33_port, B2 => n6, Y => n81);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(34), A2 => n3, B1 => 
                           data_tx_pl_34_port, B2 => n6, Y => n80);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(35), A2 => n3, B1 => 
                           data_tx_pl_35_port, B2 => n6, Y => n79);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(36), A2 => n3, B1 => 
                           data_tx_pl_36_port, B2 => n6, Y => n78);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(37), A2 => n3, B1 => 
                           data_tx_pl_37_port, B2 => n6, Y => n76);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(38), A2 => n3, B1 => 
                           data_tx_pl_38_port, B2 => n6, Y => n74);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(39), A2 => n3, B1 => 
                           data_tx_pl_39_port, B2 => n6, Y => n72);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(40), A2 => n3, B1 => 
                           data_tx_pl_40_port, B2 => n5, Y => n70);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(41), A2 => n3, B1 => 
                           data_tx_pl_41_port, B2 => n5, Y => n68);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(42), A2 => n3, B1 => 
                           data_tx_pl_42_port, B2 => n5, Y => n66);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(43), A2 => n3, B1 => 
                           data_tx_pl_43_port, B2 => n5, Y => n64);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(44), A2 => n3, B1 => 
                           data_tx_pl_44_port, B2 => n5, Y => n62);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(45), A2 => n3, B1 => 
                           data_tx_pl_45_port, B2 => n5, Y => n60);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(46), A2 => n3, B1 => 
                           data_tx_pl_46_port, B2 => n5, Y => n58);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(47), A2 => n3, B1 => 
                           data_tx_pl_47_port, B2 => n5, Y => n56);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(48), A2 => n3, B1 => 
                           data_tx_pl_48_port, B2 => n5, Y => n54);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(49), A2 => n3, B1 => 
                           data_tx_pl_49_port, B2 => n5, Y => n52);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(50), A2 => n3, B1 => 
                           data_tx_pl_50_port, B2 => n5, Y => n50);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(51), A2 => n3, B1 => 
                           data_tx_pl_51_port, B2 => n5, Y => n48);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(52), A2 => n3, B1 => 
                           data_tx_pl_52_port, B2 => n4, Y => n46);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(53), A2 => n3, B1 => 
                           data_tx_pl_53_port, B2 => n4, Y => n44);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(54), A2 => n3, B1 => 
                           data_tx_pl_54_port, B2 => n4, Y => n42);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(55), A2 => n3, B1 => 
                           data_tx_pl_55_port, B2 => n4, Y => n40);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(56), A2 => n3, B1 => 
                           data_tx_pl_56_port, B2 => n4, Y => n38);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(57), A2 => n3, B1 => 
                           data_tx_pl_57_port, B2 => n4, Y => n36);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(58), A2 => n3, B1 => 
                           data_tx_pl_58_port, B2 => n4, Y => n34);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(59), A2 => n3, B1 => 
                           data_tx_pl_59_port, B2 => n4, Y => n32);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(60), A2 => n3, B1 => 
                           data_tx_pl_60_port, B2 => n4, Y => n30);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(61), A2 => n3, B1 => 
                           data_tx_pl_61_port, B2 => n4, Y => n28);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(62), A2 => n3, B1 => 
                           data_tx_pl_62_port, B2 => n4, Y => n26);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(63), A2 => n3, B1 => 
                           data_tx_pl_63_port, B2 => n4, Y => n24);
   U68 : NAND2xp5_ASAP7_75t_R port map( A => n20, B => n22, Y => n115);
   vc_write_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n22, CLK
                           => clk, RESET => n16, SET => n1, QN => 
                           vc_write_tx_pl(0));
   vc_write_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n20, CLK
                           => clk, RESET => n16, SET => n1, QN => 
                           vc_write_tx_pl(1));
   incr_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n14, CLK => 
                           clk, RESET => n16, SET => n1, QN => incr_tx_pl(1));
   incr_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n18, CLK => 
                           clk, RESET => n16, SET => n1, QN => incr_tx_pl(0));
   data_tx_pl_reg_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n50, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_50_port);
   data_tx_pl_reg_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n52, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_49_port);
   data_tx_pl_reg_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n54, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_48_port);
   data_tx_pl_reg_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n56, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_47_port);
   data_tx_pl_reg_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n58, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_46_port);
   data_tx_pl_reg_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n60, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_45_port);
   data_tx_pl_reg_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n62, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_44_port);
   data_tx_pl_reg_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n64, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_43_port);
   data_tx_pl_reg_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n66, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_42_port);
   data_tx_pl_reg_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n68, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_41_port);
   data_tx_pl_reg_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n70, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_40_port);
   data_tx_pl_reg_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n72, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_39_port);
   data_tx_pl_reg_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n74, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_38_port);
   data_tx_pl_reg_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n76, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_37_port);
   data_tx_pl_reg_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n78, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_36_port);
   data_tx_pl_reg_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_35_port);
   data_tx_pl_reg_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n80, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_34_port);
   data_tx_pl_reg_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_33_port);
   data_tx_pl_reg_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n82, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_32_port);
   data_tx_pl_reg_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_31_port);
   data_tx_pl_reg_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n84, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_30_port);
   data_tx_pl_reg_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_9_port);
   data_tx_pl_reg_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n106, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_8_port);
   data_tx_pl_reg_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_7_port);
   data_tx_pl_reg_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n108, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_6_port);
   data_tx_pl_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_3_port);
   data_tx_pl_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n112, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_2_port);
   data_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_1_port);
   data_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n114, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_0_port);
   data_tx_pl_reg_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n24, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_63_port);
   data_tx_pl_reg_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n26, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_62_port);
   data_tx_pl_reg_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n28, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_61_port);
   data_tx_pl_reg_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n30, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_60_port);
   data_tx_pl_reg_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n32, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_59_port);
   data_tx_pl_reg_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n34, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_58_port);
   data_tx_pl_reg_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n36, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_57_port);
   data_tx_pl_reg_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n38, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_56_port);
   data_tx_pl_reg_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n40, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_55_port);
   data_tx_pl_reg_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n42, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_54_port);
   data_tx_pl_reg_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n44, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_53_port);
   data_tx_pl_reg_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n46, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_52_port);
   data_tx_pl_reg_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n48, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_51_port);
   data_tx_pl_reg_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_29_port);
   data_tx_pl_reg_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n86, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_28_port);
   data_tx_pl_reg_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_27_port);
   data_tx_pl_reg_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n88, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_26_port);
   data_tx_pl_reg_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_25_port);
   data_tx_pl_reg_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n90, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_24_port);
   data_tx_pl_reg_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_23_port);
   data_tx_pl_reg_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n92, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_22_port);
   data_tx_pl_reg_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_21_port);
   data_tx_pl_reg_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n94, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_20_port);
   data_tx_pl_reg_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_19_port);
   data_tx_pl_reg_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n96, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_18_port);
   data_tx_pl_reg_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_17_port);
   data_tx_pl_reg_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n98, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_16_port);
   data_tx_pl_reg_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_15_port);
   data_tx_pl_reg_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n100, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_14_port);
   data_tx_pl_reg_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_13_port);
   data_tx_pl_reg_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n102, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_12_port);
   data_tx_pl_reg_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_11_port);
   data_tx_pl_reg_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n104, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_10_port);
   data_tx_pl_reg_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_5_port);
   data_tx_pl_reg_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n110, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_4_port);
   U67 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U69 : INVx2_ASAP7_75t_R port map( A => rst, Y => n16);
   U70 : INVx1_ASAP7_75t_R port map( A => n12, Y => n3);
   U71 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n12);
   U72 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n10);
   U73 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n8);
   U74 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n4);
   U75 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n6);
   U76 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n5);
   U77 : INVx1_ASAP7_75t_R port map( A => incr_tx(1), Y => n14);
   U78 : INVx1_ASAP7_75t_R port map( A => incr_tx(0), Y => n18);
   U79 : INVx1_ASAP7_75t_R port map( A => vc_write_tx(1), Y => n20);
   U80 : INVx1_ASAP7_75t_R port map( A => vc_write_tx(0), Y => n22);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity output_register_vc_num2_vc_num_out2_4 is

   port( clk, rst : in std_logic;  data_tx : in std_logic_vector (63 downto 0);
         vc_write_tx, incr_tx : in std_logic_vector (1 downto 0);  data_tx_pl :
         out std_logic_vector (63 downto 0);  vc_write_tx_pl, incr_tx_pl : out 
         std_logic_vector (1 downto 0));

end output_register_vc_num2_vc_num_out2_4;

architecture SYN_rtl of output_register_vc_num2_vc_num_out2_4 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx2_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal data_tx_pl_63_port, data_tx_pl_62_port, data_tx_pl_61_port, 
      data_tx_pl_60_port, data_tx_pl_59_port, data_tx_pl_58_port, 
      data_tx_pl_57_port, data_tx_pl_56_port, data_tx_pl_55_port, 
      data_tx_pl_54_port, data_tx_pl_53_port, data_tx_pl_52_port, 
      data_tx_pl_51_port, data_tx_pl_50_port, data_tx_pl_49_port, 
      data_tx_pl_48_port, data_tx_pl_47_port, data_tx_pl_46_port, 
      data_tx_pl_45_port, data_tx_pl_44_port, data_tx_pl_43_port, 
      data_tx_pl_42_port, data_tx_pl_41_port, data_tx_pl_40_port, 
      data_tx_pl_39_port, data_tx_pl_38_port, data_tx_pl_37_port, 
      data_tx_pl_36_port, data_tx_pl_35_port, data_tx_pl_34_port, 
      data_tx_pl_33_port, data_tx_pl_32_port, data_tx_pl_31_port, 
      data_tx_pl_30_port, data_tx_pl_29_port, data_tx_pl_28_port, 
      data_tx_pl_27_port, data_tx_pl_26_port, data_tx_pl_25_port, 
      data_tx_pl_24_port, data_tx_pl_23_port, data_tx_pl_22_port, 
      data_tx_pl_21_port, data_tx_pl_20_port, data_tx_pl_19_port, 
      data_tx_pl_18_port, data_tx_pl_17_port, data_tx_pl_16_port, 
      data_tx_pl_15_port, data_tx_pl_14_port, data_tx_pl_13_port, 
      data_tx_pl_12_port, data_tx_pl_11_port, data_tx_pl_10_port, 
      data_tx_pl_9_port, data_tx_pl_8_port, data_tx_pl_7_port, 
      data_tx_pl_6_port, data_tx_pl_5_port, data_tx_pl_4_port, 
      data_tx_pl_3_port, data_tx_pl_2_port, data_tx_pl_1_port, 
      data_tx_pl_0_port, n1, n3, n4, n5, n6, n8, n10, n12, n14, n16, n18, n20, 
      n22, n24, n26, n28, n30, n32, n34, n36, n38, n40, n42, n44, n46, n48, n50
      , n52, n54, n56, n58, n60, n62, n64, n66, n68, n70, n72, n74, n76, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
      n107, n108, n109, n110, n111, n112, n113, n114, n115 : std_logic;

begin
   data_tx_pl <= ( data_tx_pl_63_port, data_tx_pl_62_port, data_tx_pl_61_port, 
      data_tx_pl_60_port, data_tx_pl_59_port, data_tx_pl_58_port, 
      data_tx_pl_57_port, data_tx_pl_56_port, data_tx_pl_55_port, 
      data_tx_pl_54_port, data_tx_pl_53_port, data_tx_pl_52_port, 
      data_tx_pl_51_port, data_tx_pl_50_port, data_tx_pl_49_port, 
      data_tx_pl_48_port, data_tx_pl_47_port, data_tx_pl_46_port, 
      data_tx_pl_45_port, data_tx_pl_44_port, data_tx_pl_43_port, 
      data_tx_pl_42_port, data_tx_pl_41_port, data_tx_pl_40_port, 
      data_tx_pl_39_port, data_tx_pl_38_port, data_tx_pl_37_port, 
      data_tx_pl_36_port, data_tx_pl_35_port, data_tx_pl_34_port, 
      data_tx_pl_33_port, data_tx_pl_32_port, data_tx_pl_31_port, 
      data_tx_pl_30_port, data_tx_pl_29_port, data_tx_pl_28_port, 
      data_tx_pl_27_port, data_tx_pl_26_port, data_tx_pl_25_port, 
      data_tx_pl_24_port, data_tx_pl_23_port, data_tx_pl_22_port, 
      data_tx_pl_21_port, data_tx_pl_20_port, data_tx_pl_19_port, 
      data_tx_pl_18_port, data_tx_pl_17_port, data_tx_pl_16_port, 
      data_tx_pl_15_port, data_tx_pl_14_port, data_tx_pl_13_port, 
      data_tx_pl_12_port, data_tx_pl_11_port, data_tx_pl_10_port, 
      data_tx_pl_9_port, data_tx_pl_8_port, data_tx_pl_7_port, 
      data_tx_pl_6_port, data_tx_pl_5_port, data_tx_pl_4_port, 
      data_tx_pl_3_port, data_tx_pl_2_port, data_tx_pl_1_port, 
      data_tx_pl_0_port );
   
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(0), A2 => n3, B1 => 
                           data_tx_pl_0_port, B2 => n12, Y => n114);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(1), A2 => n3, B1 => 
                           data_tx_pl_1_port, B2 => n12, Y => n113);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(2), A2 => n3, B1 => 
                           data_tx_pl_2_port, B2 => n12, Y => n112);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(3), A2 => n3, B1 => 
                           data_tx_pl_3_port, B2 => n12, Y => n111);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(4), A2 => n3, B1 => 
                           data_tx_pl_4_port, B2 => n10, Y => n110);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(5), A2 => n3, B1 => 
                           data_tx_pl_5_port, B2 => n10, Y => n109);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(6), A2 => n3, B1 => 
                           data_tx_pl_6_port, B2 => n10, Y => n108);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(7), A2 => n3, B1 => 
                           data_tx_pl_7_port, B2 => n10, Y => n107);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(8), A2 => n3, B1 => 
                           data_tx_pl_8_port, B2 => n10, Y => n106);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(9), A2 => n3, B1 => 
                           data_tx_pl_9_port, B2 => n10, Y => n105);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(10), A2 => n3, B1 => 
                           data_tx_pl_10_port, B2 => n10, Y => n104);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(11), A2 => n3, B1 => 
                           data_tx_pl_11_port, B2 => n10, Y => n103);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(12), A2 => n3, B1 => 
                           data_tx_pl_12_port, B2 => n10, Y => n102);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(13), A2 => n3, B1 => 
                           data_tx_pl_13_port, B2 => n10, Y => n101);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(14), A2 => n3, B1 => 
                           data_tx_pl_14_port, B2 => n10, Y => n100);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(15), A2 => n3, B1 => 
                           data_tx_pl_15_port, B2 => n10, Y => n99);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(16), A2 => n3, B1 => 
                           data_tx_pl_16_port, B2 => n8, Y => n98);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(17), A2 => n3, B1 => 
                           data_tx_pl_17_port, B2 => n8, Y => n97);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(18), A2 => n3, B1 => 
                           data_tx_pl_18_port, B2 => n8, Y => n96);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(19), A2 => n3, B1 => 
                           data_tx_pl_19_port, B2 => n8, Y => n95);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(20), A2 => n3, B1 => 
                           data_tx_pl_20_port, B2 => n8, Y => n94);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(21), A2 => n3, B1 => 
                           data_tx_pl_21_port, B2 => n8, Y => n93);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(22), A2 => n3, B1 => 
                           data_tx_pl_22_port, B2 => n8, Y => n92);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(23), A2 => n3, B1 => 
                           data_tx_pl_23_port, B2 => n8, Y => n91);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(24), A2 => n3, B1 => 
                           data_tx_pl_24_port, B2 => n8, Y => n90);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(25), A2 => n3, B1 => 
                           data_tx_pl_25_port, B2 => n8, Y => n89);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(26), A2 => n3, B1 => 
                           data_tx_pl_26_port, B2 => n8, Y => n88);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(27), A2 => n3, B1 => 
                           data_tx_pl_27_port, B2 => n8, Y => n87);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(28), A2 => n3, B1 => 
                           data_tx_pl_28_port, B2 => n6, Y => n86);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(29), A2 => n3, B1 => 
                           data_tx_pl_29_port, B2 => n6, Y => n85);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(30), A2 => n3, B1 => 
                           data_tx_pl_30_port, B2 => n6, Y => n84);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(31), A2 => n3, B1 => 
                           data_tx_pl_31_port, B2 => n6, Y => n83);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(32), A2 => n3, B1 => 
                           data_tx_pl_32_port, B2 => n6, Y => n82);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(33), A2 => n3, B1 => 
                           data_tx_pl_33_port, B2 => n6, Y => n81);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(34), A2 => n3, B1 => 
                           data_tx_pl_34_port, B2 => n6, Y => n80);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(35), A2 => n3, B1 => 
                           data_tx_pl_35_port, B2 => n6, Y => n79);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(36), A2 => n3, B1 => 
                           data_tx_pl_36_port, B2 => n6, Y => n78);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(37), A2 => n3, B1 => 
                           data_tx_pl_37_port, B2 => n6, Y => n76);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(38), A2 => n3, B1 => 
                           data_tx_pl_38_port, B2 => n6, Y => n74);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(39), A2 => n3, B1 => 
                           data_tx_pl_39_port, B2 => n6, Y => n72);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(40), A2 => n3, B1 => 
                           data_tx_pl_40_port, B2 => n5, Y => n70);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(41), A2 => n3, B1 => 
                           data_tx_pl_41_port, B2 => n5, Y => n68);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(42), A2 => n3, B1 => 
                           data_tx_pl_42_port, B2 => n5, Y => n66);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(43), A2 => n3, B1 => 
                           data_tx_pl_43_port, B2 => n5, Y => n64);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(44), A2 => n3, B1 => 
                           data_tx_pl_44_port, B2 => n5, Y => n62);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(45), A2 => n3, B1 => 
                           data_tx_pl_45_port, B2 => n5, Y => n60);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(46), A2 => n3, B1 => 
                           data_tx_pl_46_port, B2 => n5, Y => n58);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(47), A2 => n3, B1 => 
                           data_tx_pl_47_port, B2 => n5, Y => n56);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(48), A2 => n3, B1 => 
                           data_tx_pl_48_port, B2 => n5, Y => n54);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(49), A2 => n3, B1 => 
                           data_tx_pl_49_port, B2 => n5, Y => n52);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(50), A2 => n3, B1 => 
                           data_tx_pl_50_port, B2 => n5, Y => n50);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(51), A2 => n3, B1 => 
                           data_tx_pl_51_port, B2 => n5, Y => n48);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(52), A2 => n3, B1 => 
                           data_tx_pl_52_port, B2 => n4, Y => n46);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(53), A2 => n3, B1 => 
                           data_tx_pl_53_port, B2 => n4, Y => n44);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(54), A2 => n3, B1 => 
                           data_tx_pl_54_port, B2 => n4, Y => n42);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(55), A2 => n3, B1 => 
                           data_tx_pl_55_port, B2 => n4, Y => n40);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(56), A2 => n3, B1 => 
                           data_tx_pl_56_port, B2 => n4, Y => n38);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(57), A2 => n3, B1 => 
                           data_tx_pl_57_port, B2 => n4, Y => n36);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(58), A2 => n3, B1 => 
                           data_tx_pl_58_port, B2 => n4, Y => n34);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(59), A2 => n3, B1 => 
                           data_tx_pl_59_port, B2 => n4, Y => n32);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(60), A2 => n3, B1 => 
                           data_tx_pl_60_port, B2 => n4, Y => n30);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(61), A2 => n3, B1 => 
                           data_tx_pl_61_port, B2 => n4, Y => n28);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(62), A2 => n3, B1 => 
                           data_tx_pl_62_port, B2 => n4, Y => n26);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(63), A2 => n3, B1 => 
                           data_tx_pl_63_port, B2 => n4, Y => n24);
   U68 : NAND2xp5_ASAP7_75t_R port map( A => n20, B => n22, Y => n115);
   vc_write_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n20, CLK
                           => clk, RESET => n16, SET => n1, QN => 
                           vc_write_tx_pl(1));
   vc_write_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n22, CLK
                           => clk, RESET => n16, SET => n1, QN => 
                           vc_write_tx_pl(0));
   incr_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n14, CLK => 
                           clk, RESET => n16, SET => n1, QN => incr_tx_pl(1));
   incr_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n18, CLK => 
                           clk, RESET => n16, SET => n1, QN => incr_tx_pl(0));
   data_tx_pl_reg_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n50, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_50_port);
   data_tx_pl_reg_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n52, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_49_port);
   data_tx_pl_reg_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n54, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_48_port);
   data_tx_pl_reg_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n56, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_47_port);
   data_tx_pl_reg_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n58, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_46_port);
   data_tx_pl_reg_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n60, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_45_port);
   data_tx_pl_reg_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n62, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_44_port);
   data_tx_pl_reg_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n64, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_43_port);
   data_tx_pl_reg_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n66, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_42_port);
   data_tx_pl_reg_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n68, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_41_port);
   data_tx_pl_reg_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n70, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_40_port);
   data_tx_pl_reg_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n72, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_39_port);
   data_tx_pl_reg_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n74, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_38_port);
   data_tx_pl_reg_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n76, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_37_port);
   data_tx_pl_reg_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n78, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_36_port);
   data_tx_pl_reg_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_35_port);
   data_tx_pl_reg_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n80, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_34_port);
   data_tx_pl_reg_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_33_port);
   data_tx_pl_reg_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n82, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_32_port);
   data_tx_pl_reg_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_31_port);
   data_tx_pl_reg_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n84, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_30_port);
   data_tx_pl_reg_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n102, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_12_port);
   data_tx_pl_reg_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_11_port);
   data_tx_pl_reg_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n104, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_10_port);
   data_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n114, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_0_port);
   data_tx_pl_reg_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n24, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_63_port);
   data_tx_pl_reg_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n26, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_62_port);
   data_tx_pl_reg_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n28, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_61_port);
   data_tx_pl_reg_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n30, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_60_port);
   data_tx_pl_reg_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n32, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_59_port);
   data_tx_pl_reg_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n34, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_58_port);
   data_tx_pl_reg_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n36, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_57_port);
   data_tx_pl_reg_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n38, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_56_port);
   data_tx_pl_reg_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n40, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_55_port);
   data_tx_pl_reg_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n42, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_54_port);
   data_tx_pl_reg_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n44, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_53_port);
   data_tx_pl_reg_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n46, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_52_port);
   data_tx_pl_reg_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n48, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_51_port);
   data_tx_pl_reg_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_29_port);
   data_tx_pl_reg_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n86, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_28_port);
   data_tx_pl_reg_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_27_port);
   data_tx_pl_reg_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n88, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_26_port);
   data_tx_pl_reg_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_25_port);
   data_tx_pl_reg_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n90, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_24_port);
   data_tx_pl_reg_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_23_port);
   data_tx_pl_reg_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n92, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_22_port);
   data_tx_pl_reg_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_21_port);
   data_tx_pl_reg_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n94, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_20_port);
   data_tx_pl_reg_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_19_port);
   data_tx_pl_reg_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n96, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_18_port);
   data_tx_pl_reg_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_17_port);
   data_tx_pl_reg_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n98, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_16_port);
   data_tx_pl_reg_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_15_port);
   data_tx_pl_reg_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n100, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_14_port);
   data_tx_pl_reg_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_13_port);
   data_tx_pl_reg_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_9_port);
   data_tx_pl_reg_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n106, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_8_port);
   data_tx_pl_reg_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_7_port);
   data_tx_pl_reg_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n108, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_6_port);
   data_tx_pl_reg_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_5_port);
   data_tx_pl_reg_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n110, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_4_port);
   data_tx_pl_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_3_port);
   data_tx_pl_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n112, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_2_port);
   data_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_1_port);
   U67 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U69 : INVx2_ASAP7_75t_R port map( A => rst, Y => n16);
   U70 : INVx1_ASAP7_75t_R port map( A => n12, Y => n3);
   U71 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n12);
   U72 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n10);
   U73 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n8);
   U74 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n6);
   U75 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n5);
   U76 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n4);
   U77 : INVx1_ASAP7_75t_R port map( A => incr_tx(1), Y => n14);
   U78 : INVx1_ASAP7_75t_R port map( A => incr_tx(0), Y => n18);
   U79 : INVx1_ASAP7_75t_R port map( A => vc_write_tx(1), Y => n20);
   U80 : INVx1_ASAP7_75t_R port map( A => vc_write_tx(0), Y => n22);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity output_register_vc_num2_vc_num_out2_3 is

   port( clk, rst : in std_logic;  data_tx : in std_logic_vector (63 downto 0);
         vc_write_tx, incr_tx : in std_logic_vector (1 downto 0);  data_tx_pl :
         out std_logic_vector (63 downto 0);  vc_write_tx_pl, incr_tx_pl : out 
         std_logic_vector (1 downto 0));

end output_register_vc_num2_vc_num_out2_3;

architecture SYN_rtl of output_register_vc_num2_vc_num_out2_3 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx2_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal data_tx_pl_63_port, data_tx_pl_62_port, data_tx_pl_61_port, 
      data_tx_pl_60_port, data_tx_pl_59_port, data_tx_pl_58_port, 
      data_tx_pl_57_port, data_tx_pl_56_port, data_tx_pl_55_port, 
      data_tx_pl_54_port, data_tx_pl_53_port, data_tx_pl_52_port, 
      data_tx_pl_51_port, data_tx_pl_50_port, data_tx_pl_49_port, 
      data_tx_pl_48_port, data_tx_pl_47_port, data_tx_pl_46_port, 
      data_tx_pl_45_port, data_tx_pl_44_port, data_tx_pl_43_port, 
      data_tx_pl_42_port, data_tx_pl_41_port, data_tx_pl_40_port, 
      data_tx_pl_39_port, data_tx_pl_38_port, data_tx_pl_37_port, 
      data_tx_pl_36_port, data_tx_pl_35_port, data_tx_pl_34_port, 
      data_tx_pl_33_port, data_tx_pl_32_port, data_tx_pl_31_port, 
      data_tx_pl_30_port, data_tx_pl_29_port, data_tx_pl_28_port, 
      data_tx_pl_27_port, data_tx_pl_26_port, data_tx_pl_25_port, 
      data_tx_pl_24_port, data_tx_pl_23_port, data_tx_pl_22_port, 
      data_tx_pl_21_port, data_tx_pl_20_port, data_tx_pl_19_port, 
      data_tx_pl_18_port, data_tx_pl_17_port, data_tx_pl_16_port, 
      data_tx_pl_15_port, data_tx_pl_14_port, data_tx_pl_13_port, 
      data_tx_pl_12_port, data_tx_pl_11_port, data_tx_pl_10_port, 
      data_tx_pl_9_port, data_tx_pl_8_port, data_tx_pl_7_port, 
      data_tx_pl_6_port, data_tx_pl_5_port, data_tx_pl_4_port, 
      data_tx_pl_3_port, data_tx_pl_2_port, data_tx_pl_1_port, 
      data_tx_pl_0_port, n1, n3, n4, n5, n6, n8, n10, n12, n14, n16, n18, n20, 
      n22, n24, n26, n28, n30, n32, n34, n36, n38, n40, n42, n44, n46, n48, n50
      , n52, n54, n56, n58, n60, n62, n64, n66, n68, n70, n72, n74, n76, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
      n107, n108, n109, n110, n111, n112, n113, n114, n115 : std_logic;

begin
   data_tx_pl <= ( data_tx_pl_63_port, data_tx_pl_62_port, data_tx_pl_61_port, 
      data_tx_pl_60_port, data_tx_pl_59_port, data_tx_pl_58_port, 
      data_tx_pl_57_port, data_tx_pl_56_port, data_tx_pl_55_port, 
      data_tx_pl_54_port, data_tx_pl_53_port, data_tx_pl_52_port, 
      data_tx_pl_51_port, data_tx_pl_50_port, data_tx_pl_49_port, 
      data_tx_pl_48_port, data_tx_pl_47_port, data_tx_pl_46_port, 
      data_tx_pl_45_port, data_tx_pl_44_port, data_tx_pl_43_port, 
      data_tx_pl_42_port, data_tx_pl_41_port, data_tx_pl_40_port, 
      data_tx_pl_39_port, data_tx_pl_38_port, data_tx_pl_37_port, 
      data_tx_pl_36_port, data_tx_pl_35_port, data_tx_pl_34_port, 
      data_tx_pl_33_port, data_tx_pl_32_port, data_tx_pl_31_port, 
      data_tx_pl_30_port, data_tx_pl_29_port, data_tx_pl_28_port, 
      data_tx_pl_27_port, data_tx_pl_26_port, data_tx_pl_25_port, 
      data_tx_pl_24_port, data_tx_pl_23_port, data_tx_pl_22_port, 
      data_tx_pl_21_port, data_tx_pl_20_port, data_tx_pl_19_port, 
      data_tx_pl_18_port, data_tx_pl_17_port, data_tx_pl_16_port, 
      data_tx_pl_15_port, data_tx_pl_14_port, data_tx_pl_13_port, 
      data_tx_pl_12_port, data_tx_pl_11_port, data_tx_pl_10_port, 
      data_tx_pl_9_port, data_tx_pl_8_port, data_tx_pl_7_port, 
      data_tx_pl_6_port, data_tx_pl_5_port, data_tx_pl_4_port, 
      data_tx_pl_3_port, data_tx_pl_2_port, data_tx_pl_1_port, 
      data_tx_pl_0_port );
   
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(0), A2 => n3, B1 => 
                           data_tx_pl_0_port, B2 => n12, Y => n114);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(1), A2 => n3, B1 => 
                           data_tx_pl_1_port, B2 => n12, Y => n113);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(2), A2 => n3, B1 => 
                           data_tx_pl_2_port, B2 => n12, Y => n112);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(3), A2 => n3, B1 => 
                           data_tx_pl_3_port, B2 => n12, Y => n111);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(4), A2 => n3, B1 => 
                           data_tx_pl_4_port, B2 => n10, Y => n110);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(5), A2 => n3, B1 => 
                           data_tx_pl_5_port, B2 => n10, Y => n109);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(6), A2 => n3, B1 => 
                           data_tx_pl_6_port, B2 => n10, Y => n108);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(7), A2 => n3, B1 => 
                           data_tx_pl_7_port, B2 => n10, Y => n107);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(8), A2 => n3, B1 => 
                           data_tx_pl_8_port, B2 => n10, Y => n106);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(9), A2 => n3, B1 => 
                           data_tx_pl_9_port, B2 => n10, Y => n105);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(10), A2 => n3, B1 => 
                           data_tx_pl_10_port, B2 => n10, Y => n104);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(11), A2 => n3, B1 => 
                           data_tx_pl_11_port, B2 => n10, Y => n103);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(12), A2 => n3, B1 => 
                           data_tx_pl_12_port, B2 => n10, Y => n102);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(13), A2 => n3, B1 => 
                           data_tx_pl_13_port, B2 => n10, Y => n101);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(14), A2 => n3, B1 => 
                           data_tx_pl_14_port, B2 => n10, Y => n100);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(15), A2 => n3, B1 => 
                           data_tx_pl_15_port, B2 => n10, Y => n99);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(16), A2 => n3, B1 => 
                           data_tx_pl_16_port, B2 => n8, Y => n98);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(17), A2 => n3, B1 => 
                           data_tx_pl_17_port, B2 => n8, Y => n97);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(18), A2 => n3, B1 => 
                           data_tx_pl_18_port, B2 => n8, Y => n96);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(19), A2 => n3, B1 => 
                           data_tx_pl_19_port, B2 => n8, Y => n95);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(20), A2 => n3, B1 => 
                           data_tx_pl_20_port, B2 => n8, Y => n94);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(21), A2 => n3, B1 => 
                           data_tx_pl_21_port, B2 => n8, Y => n93);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(22), A2 => n3, B1 => 
                           data_tx_pl_22_port, B2 => n8, Y => n92);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(23), A2 => n3, B1 => 
                           data_tx_pl_23_port, B2 => n8, Y => n91);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(24), A2 => n3, B1 => 
                           data_tx_pl_24_port, B2 => n8, Y => n90);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(25), A2 => n3, B1 => 
                           data_tx_pl_25_port, B2 => n8, Y => n89);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(26), A2 => n3, B1 => 
                           data_tx_pl_26_port, B2 => n8, Y => n88);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(27), A2 => n3, B1 => 
                           data_tx_pl_27_port, B2 => n8, Y => n87);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(28), A2 => n3, B1 => 
                           data_tx_pl_28_port, B2 => n6, Y => n86);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(29), A2 => n3, B1 => 
                           data_tx_pl_29_port, B2 => n6, Y => n85);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(30), A2 => n3, B1 => 
                           data_tx_pl_30_port, B2 => n6, Y => n84);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(31), A2 => n3, B1 => 
                           data_tx_pl_31_port, B2 => n6, Y => n83);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(32), A2 => n3, B1 => 
                           data_tx_pl_32_port, B2 => n6, Y => n82);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(33), A2 => n3, B1 => 
                           data_tx_pl_33_port, B2 => n6, Y => n81);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(34), A2 => n3, B1 => 
                           data_tx_pl_34_port, B2 => n6, Y => n80);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(35), A2 => n3, B1 => 
                           data_tx_pl_35_port, B2 => n6, Y => n79);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(36), A2 => n3, B1 => 
                           data_tx_pl_36_port, B2 => n6, Y => n78);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(37), A2 => n3, B1 => 
                           data_tx_pl_37_port, B2 => n6, Y => n76);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(38), A2 => n3, B1 => 
                           data_tx_pl_38_port, B2 => n6, Y => n74);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(39), A2 => n3, B1 => 
                           data_tx_pl_39_port, B2 => n6, Y => n72);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(40), A2 => n3, B1 => 
                           data_tx_pl_40_port, B2 => n5, Y => n70);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(41), A2 => n3, B1 => 
                           data_tx_pl_41_port, B2 => n5, Y => n68);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(42), A2 => n3, B1 => 
                           data_tx_pl_42_port, B2 => n5, Y => n66);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(43), A2 => n3, B1 => 
                           data_tx_pl_43_port, B2 => n5, Y => n64);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(44), A2 => n3, B1 => 
                           data_tx_pl_44_port, B2 => n5, Y => n62);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(45), A2 => n3, B1 => 
                           data_tx_pl_45_port, B2 => n5, Y => n60);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(46), A2 => n3, B1 => 
                           data_tx_pl_46_port, B2 => n5, Y => n58);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(47), A2 => n3, B1 => 
                           data_tx_pl_47_port, B2 => n5, Y => n56);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(48), A2 => n3, B1 => 
                           data_tx_pl_48_port, B2 => n5, Y => n54);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(49), A2 => n3, B1 => 
                           data_tx_pl_49_port, B2 => n5, Y => n52);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(50), A2 => n3, B1 => 
                           data_tx_pl_50_port, B2 => n5, Y => n50);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(51), A2 => n3, B1 => 
                           data_tx_pl_51_port, B2 => n5, Y => n48);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(52), A2 => n3, B1 => 
                           data_tx_pl_52_port, B2 => n4, Y => n46);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(53), A2 => n3, B1 => 
                           data_tx_pl_53_port, B2 => n4, Y => n44);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(54), A2 => n3, B1 => 
                           data_tx_pl_54_port, B2 => n4, Y => n42);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(55), A2 => n3, B1 => 
                           data_tx_pl_55_port, B2 => n4, Y => n40);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(56), A2 => n3, B1 => 
                           data_tx_pl_56_port, B2 => n4, Y => n38);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(57), A2 => n3, B1 => 
                           data_tx_pl_57_port, B2 => n4, Y => n36);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(58), A2 => n3, B1 => 
                           data_tx_pl_58_port, B2 => n4, Y => n34);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(59), A2 => n3, B1 => 
                           data_tx_pl_59_port, B2 => n4, Y => n32);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(60), A2 => n3, B1 => 
                           data_tx_pl_60_port, B2 => n4, Y => n30);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(61), A2 => n3, B1 => 
                           data_tx_pl_61_port, B2 => n4, Y => n28);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(62), A2 => n3, B1 => 
                           data_tx_pl_62_port, B2 => n4, Y => n26);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(63), A2 => n3, B1 => 
                           data_tx_pl_63_port, B2 => n4, Y => n24);
   U68 : NAND2xp5_ASAP7_75t_R port map( A => n20, B => n22, Y => n115);
   vc_write_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n22, CLK
                           => clk, RESET => n16, SET => n1, QN => 
                           vc_write_tx_pl(0));
   vc_write_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n20, CLK
                           => clk, RESET => n16, SET => n1, QN => 
                           vc_write_tx_pl(1));
   incr_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n14, CLK => 
                           clk, RESET => n16, SET => n1, QN => incr_tx_pl(1));
   incr_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n18, CLK => 
                           clk, RESET => n16, SET => n1, QN => incr_tx_pl(0));
   data_tx_pl_reg_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n50, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_50_port);
   data_tx_pl_reg_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n52, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_49_port);
   data_tx_pl_reg_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n54, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_48_port);
   data_tx_pl_reg_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n56, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_47_port);
   data_tx_pl_reg_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n58, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_46_port);
   data_tx_pl_reg_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n60, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_45_port);
   data_tx_pl_reg_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n62, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_44_port);
   data_tx_pl_reg_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n64, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_43_port);
   data_tx_pl_reg_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n66, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_42_port);
   data_tx_pl_reg_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n68, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_41_port);
   data_tx_pl_reg_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n70, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_40_port);
   data_tx_pl_reg_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n72, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_39_port);
   data_tx_pl_reg_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n74, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_38_port);
   data_tx_pl_reg_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n76, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_37_port);
   data_tx_pl_reg_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n78, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_36_port);
   data_tx_pl_reg_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_35_port);
   data_tx_pl_reg_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n80, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_34_port);
   data_tx_pl_reg_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_33_port);
   data_tx_pl_reg_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n82, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_32_port);
   data_tx_pl_reg_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_31_port);
   data_tx_pl_reg_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n84, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_30_port);
   data_tx_pl_reg_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_9_port);
   data_tx_pl_reg_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n106, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_8_port);
   data_tx_pl_reg_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_7_port);
   data_tx_pl_reg_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n108, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_6_port);
   data_tx_pl_reg_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n24, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_63_port);
   data_tx_pl_reg_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n26, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_62_port);
   data_tx_pl_reg_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n28, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_61_port);
   data_tx_pl_reg_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n30, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_60_port);
   data_tx_pl_reg_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n32, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_59_port);
   data_tx_pl_reg_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n34, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_58_port);
   data_tx_pl_reg_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n36, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_57_port);
   data_tx_pl_reg_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n38, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_56_port);
   data_tx_pl_reg_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n40, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_55_port);
   data_tx_pl_reg_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n42, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_54_port);
   data_tx_pl_reg_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n44, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_53_port);
   data_tx_pl_reg_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n46, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_52_port);
   data_tx_pl_reg_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n48, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_51_port);
   data_tx_pl_reg_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_29_port);
   data_tx_pl_reg_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n86, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_28_port);
   data_tx_pl_reg_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_27_port);
   data_tx_pl_reg_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n88, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_26_port);
   data_tx_pl_reg_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_25_port);
   data_tx_pl_reg_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n90, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_24_port);
   data_tx_pl_reg_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_23_port);
   data_tx_pl_reg_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n92, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_22_port);
   data_tx_pl_reg_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_21_port);
   data_tx_pl_reg_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n94, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_20_port);
   data_tx_pl_reg_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_19_port);
   data_tx_pl_reg_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n96, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_18_port);
   data_tx_pl_reg_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_17_port);
   data_tx_pl_reg_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n98, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_16_port);
   data_tx_pl_reg_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_15_port);
   data_tx_pl_reg_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n100, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_14_port);
   data_tx_pl_reg_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_13_port);
   data_tx_pl_reg_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n102, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_12_port);
   data_tx_pl_reg_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_11_port);
   data_tx_pl_reg_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n104, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_10_port);
   data_tx_pl_reg_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_5_port);
   data_tx_pl_reg_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n110, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_4_port);
   data_tx_pl_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_3_port);
   data_tx_pl_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n112, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_2_port);
   data_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_1_port);
   data_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n114, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_0_port);
   U67 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U69 : INVx2_ASAP7_75t_R port map( A => rst, Y => n16);
   U70 : INVx1_ASAP7_75t_R port map( A => n12, Y => n3);
   U71 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n12);
   U72 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n10);
   U73 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n8);
   U74 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n6);
   U75 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n5);
   U76 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n4);
   U77 : INVx1_ASAP7_75t_R port map( A => incr_tx(1), Y => n14);
   U78 : INVx1_ASAP7_75t_R port map( A => incr_tx(0), Y => n18);
   U79 : INVx1_ASAP7_75t_R port map( A => vc_write_tx(1), Y => n20);
   U80 : INVx1_ASAP7_75t_R port map( A => vc_write_tx(0), Y => n22);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity output_register_vc_num2_vc_num_out2_2 is

   port( clk, rst : in std_logic;  data_tx : in std_logic_vector (63 downto 0);
         vc_write_tx, incr_tx : in std_logic_vector (1 downto 0);  data_tx_pl :
         out std_logic_vector (63 downto 0);  vc_write_tx_pl, incr_tx_pl : out 
         std_logic_vector (1 downto 0));

end output_register_vc_num2_vc_num_out2_2;

architecture SYN_rtl of output_register_vc_num2_vc_num_out2_2 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx2_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal data_tx_pl_63_port, data_tx_pl_62_port, data_tx_pl_61_port, 
      data_tx_pl_60_port, data_tx_pl_59_port, data_tx_pl_58_port, 
      data_tx_pl_57_port, data_tx_pl_56_port, data_tx_pl_55_port, 
      data_tx_pl_54_port, data_tx_pl_53_port, data_tx_pl_52_port, 
      data_tx_pl_51_port, data_tx_pl_50_port, data_tx_pl_49_port, 
      data_tx_pl_48_port, data_tx_pl_47_port, data_tx_pl_46_port, 
      data_tx_pl_45_port, data_tx_pl_44_port, data_tx_pl_43_port, 
      data_tx_pl_42_port, data_tx_pl_41_port, data_tx_pl_40_port, 
      data_tx_pl_39_port, data_tx_pl_38_port, data_tx_pl_37_port, 
      data_tx_pl_36_port, data_tx_pl_35_port, data_tx_pl_34_port, 
      data_tx_pl_33_port, data_tx_pl_32_port, data_tx_pl_31_port, 
      data_tx_pl_30_port, data_tx_pl_29_port, data_tx_pl_28_port, 
      data_tx_pl_27_port, data_tx_pl_26_port, data_tx_pl_25_port, 
      data_tx_pl_24_port, data_tx_pl_23_port, data_tx_pl_22_port, 
      data_tx_pl_21_port, data_tx_pl_20_port, data_tx_pl_19_port, 
      data_tx_pl_18_port, data_tx_pl_17_port, data_tx_pl_16_port, 
      data_tx_pl_15_port, data_tx_pl_14_port, data_tx_pl_13_port, 
      data_tx_pl_12_port, data_tx_pl_11_port, data_tx_pl_10_port, 
      data_tx_pl_9_port, data_tx_pl_8_port, data_tx_pl_7_port, 
      data_tx_pl_6_port, data_tx_pl_5_port, data_tx_pl_4_port, 
      data_tx_pl_3_port, data_tx_pl_2_port, data_tx_pl_1_port, 
      data_tx_pl_0_port, n1, n3, n4, n5, n6, n8, n10, n12, n14, n16, n18, n20, 
      n22, n24, n26, n28, n30, n32, n34, n36, n38, n40, n42, n44, n46, n48, n50
      , n52, n54, n56, n58, n60, n62, n64, n66, n68, n70, n72, n74, n76, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
      n107, n108, n109, n110, n111, n112, n113, n114, n115 : std_logic;

begin
   data_tx_pl <= ( data_tx_pl_63_port, data_tx_pl_62_port, data_tx_pl_61_port, 
      data_tx_pl_60_port, data_tx_pl_59_port, data_tx_pl_58_port, 
      data_tx_pl_57_port, data_tx_pl_56_port, data_tx_pl_55_port, 
      data_tx_pl_54_port, data_tx_pl_53_port, data_tx_pl_52_port, 
      data_tx_pl_51_port, data_tx_pl_50_port, data_tx_pl_49_port, 
      data_tx_pl_48_port, data_tx_pl_47_port, data_tx_pl_46_port, 
      data_tx_pl_45_port, data_tx_pl_44_port, data_tx_pl_43_port, 
      data_tx_pl_42_port, data_tx_pl_41_port, data_tx_pl_40_port, 
      data_tx_pl_39_port, data_tx_pl_38_port, data_tx_pl_37_port, 
      data_tx_pl_36_port, data_tx_pl_35_port, data_tx_pl_34_port, 
      data_tx_pl_33_port, data_tx_pl_32_port, data_tx_pl_31_port, 
      data_tx_pl_30_port, data_tx_pl_29_port, data_tx_pl_28_port, 
      data_tx_pl_27_port, data_tx_pl_26_port, data_tx_pl_25_port, 
      data_tx_pl_24_port, data_tx_pl_23_port, data_tx_pl_22_port, 
      data_tx_pl_21_port, data_tx_pl_20_port, data_tx_pl_19_port, 
      data_tx_pl_18_port, data_tx_pl_17_port, data_tx_pl_16_port, 
      data_tx_pl_15_port, data_tx_pl_14_port, data_tx_pl_13_port, 
      data_tx_pl_12_port, data_tx_pl_11_port, data_tx_pl_10_port, 
      data_tx_pl_9_port, data_tx_pl_8_port, data_tx_pl_7_port, 
      data_tx_pl_6_port, data_tx_pl_5_port, data_tx_pl_4_port, 
      data_tx_pl_3_port, data_tx_pl_2_port, data_tx_pl_1_port, 
      data_tx_pl_0_port );
   
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(0), A2 => n3, B1 => 
                           data_tx_pl_0_port, B2 => n12, Y => n114);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(1), A2 => n3, B1 => 
                           data_tx_pl_1_port, B2 => n12, Y => n113);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(2), A2 => n3, B1 => 
                           data_tx_pl_2_port, B2 => n12, Y => n112);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(3), A2 => n3, B1 => 
                           data_tx_pl_3_port, B2 => n12, Y => n111);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(4), A2 => n3, B1 => 
                           data_tx_pl_4_port, B2 => n10, Y => n110);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(5), A2 => n3, B1 => 
                           data_tx_pl_5_port, B2 => n10, Y => n109);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(6), A2 => n3, B1 => 
                           data_tx_pl_6_port, B2 => n10, Y => n108);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(7), A2 => n3, B1 => 
                           data_tx_pl_7_port, B2 => n10, Y => n107);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(8), A2 => n3, B1 => 
                           data_tx_pl_8_port, B2 => n10, Y => n106);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(9), A2 => n3, B1 => 
                           data_tx_pl_9_port, B2 => n10, Y => n105);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(10), A2 => n3, B1 => 
                           data_tx_pl_10_port, B2 => n10, Y => n104);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(11), A2 => n3, B1 => 
                           data_tx_pl_11_port, B2 => n10, Y => n103);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(12), A2 => n3, B1 => 
                           data_tx_pl_12_port, B2 => n10, Y => n102);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(13), A2 => n3, B1 => 
                           data_tx_pl_13_port, B2 => n10, Y => n101);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(14), A2 => n3, B1 => 
                           data_tx_pl_14_port, B2 => n10, Y => n100);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(15), A2 => n3, B1 => 
                           data_tx_pl_15_port, B2 => n10, Y => n99);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(16), A2 => n3, B1 => 
                           data_tx_pl_16_port, B2 => n8, Y => n98);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(17), A2 => n3, B1 => 
                           data_tx_pl_17_port, B2 => n8, Y => n97);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(18), A2 => n3, B1 => 
                           data_tx_pl_18_port, B2 => n8, Y => n96);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(19), A2 => n3, B1 => 
                           data_tx_pl_19_port, B2 => n8, Y => n95);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(20), A2 => n3, B1 => 
                           data_tx_pl_20_port, B2 => n8, Y => n94);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(21), A2 => n3, B1 => 
                           data_tx_pl_21_port, B2 => n8, Y => n93);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(22), A2 => n3, B1 => 
                           data_tx_pl_22_port, B2 => n8, Y => n92);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(23), A2 => n3, B1 => 
                           data_tx_pl_23_port, B2 => n8, Y => n91);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(24), A2 => n3, B1 => 
                           data_tx_pl_24_port, B2 => n8, Y => n90);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(25), A2 => n3, B1 => 
                           data_tx_pl_25_port, B2 => n8, Y => n89);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(26), A2 => n3, B1 => 
                           data_tx_pl_26_port, B2 => n8, Y => n88);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(27), A2 => n3, B1 => 
                           data_tx_pl_27_port, B2 => n8, Y => n87);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(28), A2 => n3, B1 => 
                           data_tx_pl_28_port, B2 => n6, Y => n86);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(29), A2 => n3, B1 => 
                           data_tx_pl_29_port, B2 => n6, Y => n85);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(30), A2 => n3, B1 => 
                           data_tx_pl_30_port, B2 => n6, Y => n84);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(31), A2 => n3, B1 => 
                           data_tx_pl_31_port, B2 => n6, Y => n83);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(32), A2 => n3, B1 => 
                           data_tx_pl_32_port, B2 => n6, Y => n82);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(33), A2 => n3, B1 => 
                           data_tx_pl_33_port, B2 => n6, Y => n81);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(34), A2 => n3, B1 => 
                           data_tx_pl_34_port, B2 => n6, Y => n80);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(35), A2 => n3, B1 => 
                           data_tx_pl_35_port, B2 => n6, Y => n79);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(36), A2 => n3, B1 => 
                           data_tx_pl_36_port, B2 => n6, Y => n78);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(37), A2 => n3, B1 => 
                           data_tx_pl_37_port, B2 => n6, Y => n76);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(38), A2 => n3, B1 => 
                           data_tx_pl_38_port, B2 => n6, Y => n74);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(39), A2 => n3, B1 => 
                           data_tx_pl_39_port, B2 => n6, Y => n72);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(40), A2 => n3, B1 => 
                           data_tx_pl_40_port, B2 => n5, Y => n70);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(41), A2 => n3, B1 => 
                           data_tx_pl_41_port, B2 => n5, Y => n68);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(42), A2 => n3, B1 => 
                           data_tx_pl_42_port, B2 => n5, Y => n66);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(43), A2 => n3, B1 => 
                           data_tx_pl_43_port, B2 => n5, Y => n64);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(44), A2 => n3, B1 => 
                           data_tx_pl_44_port, B2 => n5, Y => n62);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(45), A2 => n3, B1 => 
                           data_tx_pl_45_port, B2 => n5, Y => n60);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(46), A2 => n3, B1 => 
                           data_tx_pl_46_port, B2 => n5, Y => n58);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(47), A2 => n3, B1 => 
                           data_tx_pl_47_port, B2 => n5, Y => n56);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(48), A2 => n3, B1 => 
                           data_tx_pl_48_port, B2 => n5, Y => n54);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(49), A2 => n3, B1 => 
                           data_tx_pl_49_port, B2 => n5, Y => n52);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(50), A2 => n3, B1 => 
                           data_tx_pl_50_port, B2 => n5, Y => n50);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(51), A2 => n3, B1 => 
                           data_tx_pl_51_port, B2 => n5, Y => n48);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(52), A2 => n3, B1 => 
                           data_tx_pl_52_port, B2 => n4, Y => n46);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(53), A2 => n3, B1 => 
                           data_tx_pl_53_port, B2 => n4, Y => n44);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(54), A2 => n3, B1 => 
                           data_tx_pl_54_port, B2 => n4, Y => n42);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(55), A2 => n3, B1 => 
                           data_tx_pl_55_port, B2 => n4, Y => n40);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(56), A2 => n3, B1 => 
                           data_tx_pl_56_port, B2 => n4, Y => n38);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(57), A2 => n3, B1 => 
                           data_tx_pl_57_port, B2 => n4, Y => n36);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(58), A2 => n3, B1 => 
                           data_tx_pl_58_port, B2 => n4, Y => n34);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(59), A2 => n3, B1 => 
                           data_tx_pl_59_port, B2 => n4, Y => n32);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(60), A2 => n3, B1 => 
                           data_tx_pl_60_port, B2 => n4, Y => n30);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(61), A2 => n3, B1 => 
                           data_tx_pl_61_port, B2 => n4, Y => n28);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(62), A2 => n3, B1 => 
                           data_tx_pl_62_port, B2 => n4, Y => n26);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(63), A2 => n3, B1 => 
                           data_tx_pl_63_port, B2 => n4, Y => n24);
   U68 : NAND2xp5_ASAP7_75t_R port map( A => n20, B => n22, Y => n115);
   vc_write_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n22, CLK
                           => clk, RESET => n16, SET => n1, QN => 
                           vc_write_tx_pl(0));
   vc_write_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n20, CLK
                           => clk, RESET => n16, SET => n1, QN => 
                           vc_write_tx_pl(1));
   incr_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n14, CLK => 
                           clk, RESET => n16, SET => n1, QN => incr_tx_pl(1));
   incr_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n18, CLK => 
                           clk, RESET => n16, SET => n1, QN => incr_tx_pl(0));
   data_tx_pl_reg_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n50, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_50_port);
   data_tx_pl_reg_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n52, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_49_port);
   data_tx_pl_reg_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n54, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_48_port);
   data_tx_pl_reg_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n56, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_47_port);
   data_tx_pl_reg_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n58, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_46_port);
   data_tx_pl_reg_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n60, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_45_port);
   data_tx_pl_reg_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n62, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_44_port);
   data_tx_pl_reg_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n64, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_43_port);
   data_tx_pl_reg_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n66, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_42_port);
   data_tx_pl_reg_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n68, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_41_port);
   data_tx_pl_reg_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n70, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_40_port);
   data_tx_pl_reg_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n72, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_39_port);
   data_tx_pl_reg_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n74, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_38_port);
   data_tx_pl_reg_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n76, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_37_port);
   data_tx_pl_reg_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n78, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_36_port);
   data_tx_pl_reg_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_35_port);
   data_tx_pl_reg_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n80, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_34_port);
   data_tx_pl_reg_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_33_port);
   data_tx_pl_reg_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n82, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_32_port);
   data_tx_pl_reg_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_31_port);
   data_tx_pl_reg_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n84, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_30_port);
   data_tx_pl_reg_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_19_port);
   data_tx_pl_reg_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n96, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_18_port);
   data_tx_pl_reg_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_17_port);
   data_tx_pl_reg_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n98, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_16_port);
   data_tx_pl_reg_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_15_port);
   data_tx_pl_reg_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n100, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_14_port);
   data_tx_pl_reg_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_13_port);
   data_tx_pl_reg_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n102, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_12_port);
   data_tx_pl_reg_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_11_port);
   data_tx_pl_reg_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n104, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_10_port);
   data_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_1_port);
   data_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n114, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_0_port);
   data_tx_pl_reg_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n24, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_63_port);
   data_tx_pl_reg_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n26, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_62_port);
   data_tx_pl_reg_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n28, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_61_port);
   data_tx_pl_reg_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n30, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_60_port);
   data_tx_pl_reg_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n32, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_59_port);
   data_tx_pl_reg_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n34, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_58_port);
   data_tx_pl_reg_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n36, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_57_port);
   data_tx_pl_reg_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_9_port);
   data_tx_pl_reg_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n106, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_8_port);
   data_tx_pl_reg_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_7_port);
   data_tx_pl_reg_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n108, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_6_port);
   data_tx_pl_reg_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_5_port);
   data_tx_pl_reg_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n38, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_56_port);
   data_tx_pl_reg_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n40, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_55_port);
   data_tx_pl_reg_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n42, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_54_port);
   data_tx_pl_reg_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n44, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_53_port);
   data_tx_pl_reg_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n46, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_52_port);
   data_tx_pl_reg_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n48, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_51_port);
   data_tx_pl_reg_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_29_port);
   data_tx_pl_reg_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n86, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_28_port);
   data_tx_pl_reg_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_27_port);
   data_tx_pl_reg_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n88, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_26_port);
   data_tx_pl_reg_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_25_port);
   data_tx_pl_reg_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n90, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_24_port);
   data_tx_pl_reg_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_23_port);
   data_tx_pl_reg_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n92, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_22_port);
   data_tx_pl_reg_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_21_port);
   data_tx_pl_reg_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n94, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_20_port);
   data_tx_pl_reg_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n110, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_4_port);
   data_tx_pl_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_3_port);
   data_tx_pl_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n112, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_2_port);
   U67 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U69 : INVx2_ASAP7_75t_R port map( A => rst, Y => n16);
   U70 : INVx1_ASAP7_75t_R port map( A => n12, Y => n3);
   U71 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n12);
   U72 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n10);
   U73 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n8);
   U74 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n4);
   U75 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n6);
   U76 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n5);
   U77 : INVx1_ASAP7_75t_R port map( A => incr_tx(1), Y => n14);
   U78 : INVx1_ASAP7_75t_R port map( A => incr_tx(0), Y => n18);
   U79 : INVx1_ASAP7_75t_R port map( A => vc_write_tx(1), Y => n20);
   U80 : INVx1_ASAP7_75t_R port map( A => vc_write_tx(0), Y => n22);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity output_register_vc_num2_vc_num_out2_1 is

   port( clk, rst : in std_logic;  data_tx : in std_logic_vector (63 downto 0);
         vc_write_tx, incr_tx : in std_logic_vector (1 downto 0);  data_tx_pl :
         out std_logic_vector (63 downto 0);  vc_write_tx_pl, incr_tx_pl : out 
         std_logic_vector (1 downto 0));

end output_register_vc_num2_vc_num_out2_1;

architecture SYN_rtl of output_register_vc_num2_vc_num_out2_1 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx2_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal data_tx_pl_63_port, data_tx_pl_62_port, data_tx_pl_61_port, 
      data_tx_pl_60_port, data_tx_pl_59_port, data_tx_pl_58_port, 
      data_tx_pl_57_port, data_tx_pl_56_port, data_tx_pl_55_port, 
      data_tx_pl_54_port, data_tx_pl_53_port, data_tx_pl_52_port, 
      data_tx_pl_51_port, data_tx_pl_50_port, data_tx_pl_49_port, 
      data_tx_pl_48_port, data_tx_pl_47_port, data_tx_pl_46_port, 
      data_tx_pl_45_port, data_tx_pl_44_port, data_tx_pl_43_port, 
      data_tx_pl_42_port, data_tx_pl_41_port, data_tx_pl_40_port, 
      data_tx_pl_39_port, data_tx_pl_38_port, data_tx_pl_37_port, 
      data_tx_pl_36_port, data_tx_pl_35_port, data_tx_pl_34_port, 
      data_tx_pl_33_port, data_tx_pl_32_port, data_tx_pl_31_port, 
      data_tx_pl_30_port, data_tx_pl_29_port, data_tx_pl_28_port, 
      data_tx_pl_27_port, data_tx_pl_26_port, data_tx_pl_25_port, 
      data_tx_pl_24_port, data_tx_pl_23_port, data_tx_pl_22_port, 
      data_tx_pl_21_port, data_tx_pl_20_port, data_tx_pl_19_port, 
      data_tx_pl_18_port, data_tx_pl_17_port, data_tx_pl_16_port, 
      data_tx_pl_15_port, data_tx_pl_14_port, data_tx_pl_13_port, 
      data_tx_pl_12_port, data_tx_pl_11_port, data_tx_pl_10_port, 
      data_tx_pl_9_port, data_tx_pl_8_port, data_tx_pl_7_port, 
      data_tx_pl_6_port, data_tx_pl_5_port, data_tx_pl_4_port, 
      data_tx_pl_3_port, data_tx_pl_2_port, data_tx_pl_1_port, 
      data_tx_pl_0_port, n1, n3, n4, n5, n6, n8, n10, n12, n14, n16, n18, n20, 
      n22, n24, n26, n28, n30, n32, n34, n36, n38, n40, n42, n44, n46, n48, n50
      , n52, n54, n56, n58, n60, n62, n64, n66, n68, n70, n72, n74, n76, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
      n107, n108, n109, n110, n111, n112, n113, n114, n115 : std_logic;

begin
   data_tx_pl <= ( data_tx_pl_63_port, data_tx_pl_62_port, data_tx_pl_61_port, 
      data_tx_pl_60_port, data_tx_pl_59_port, data_tx_pl_58_port, 
      data_tx_pl_57_port, data_tx_pl_56_port, data_tx_pl_55_port, 
      data_tx_pl_54_port, data_tx_pl_53_port, data_tx_pl_52_port, 
      data_tx_pl_51_port, data_tx_pl_50_port, data_tx_pl_49_port, 
      data_tx_pl_48_port, data_tx_pl_47_port, data_tx_pl_46_port, 
      data_tx_pl_45_port, data_tx_pl_44_port, data_tx_pl_43_port, 
      data_tx_pl_42_port, data_tx_pl_41_port, data_tx_pl_40_port, 
      data_tx_pl_39_port, data_tx_pl_38_port, data_tx_pl_37_port, 
      data_tx_pl_36_port, data_tx_pl_35_port, data_tx_pl_34_port, 
      data_tx_pl_33_port, data_tx_pl_32_port, data_tx_pl_31_port, 
      data_tx_pl_30_port, data_tx_pl_29_port, data_tx_pl_28_port, 
      data_tx_pl_27_port, data_tx_pl_26_port, data_tx_pl_25_port, 
      data_tx_pl_24_port, data_tx_pl_23_port, data_tx_pl_22_port, 
      data_tx_pl_21_port, data_tx_pl_20_port, data_tx_pl_19_port, 
      data_tx_pl_18_port, data_tx_pl_17_port, data_tx_pl_16_port, 
      data_tx_pl_15_port, data_tx_pl_14_port, data_tx_pl_13_port, 
      data_tx_pl_12_port, data_tx_pl_11_port, data_tx_pl_10_port, 
      data_tx_pl_9_port, data_tx_pl_8_port, data_tx_pl_7_port, 
      data_tx_pl_6_port, data_tx_pl_5_port, data_tx_pl_4_port, 
      data_tx_pl_3_port, data_tx_pl_2_port, data_tx_pl_1_port, 
      data_tx_pl_0_port );
   
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(0), A2 => n3, B1 => 
                           data_tx_pl_0_port, B2 => n12, Y => n114);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(1), A2 => n3, B1 => 
                           data_tx_pl_1_port, B2 => n12, Y => n113);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(2), A2 => n3, B1 => 
                           data_tx_pl_2_port, B2 => n12, Y => n112);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(3), A2 => n3, B1 => 
                           data_tx_pl_3_port, B2 => n12, Y => n111);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(4), A2 => n3, B1 => 
                           data_tx_pl_4_port, B2 => n10, Y => n110);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(5), A2 => n3, B1 => 
                           data_tx_pl_5_port, B2 => n10, Y => n109);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(6), A2 => n3, B1 => 
                           data_tx_pl_6_port, B2 => n10, Y => n108);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(7), A2 => n3, B1 => 
                           data_tx_pl_7_port, B2 => n10, Y => n107);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(8), A2 => n3, B1 => 
                           data_tx_pl_8_port, B2 => n10, Y => n106);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(9), A2 => n3, B1 => 
                           data_tx_pl_9_port, B2 => n10, Y => n105);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(10), A2 => n3, B1 => 
                           data_tx_pl_10_port, B2 => n10, Y => n104);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(11), A2 => n3, B1 => 
                           data_tx_pl_11_port, B2 => n10, Y => n103);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(12), A2 => n3, B1 => 
                           data_tx_pl_12_port, B2 => n10, Y => n102);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(13), A2 => n3, B1 => 
                           data_tx_pl_13_port, B2 => n10, Y => n101);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(14), A2 => n3, B1 => 
                           data_tx_pl_14_port, B2 => n10, Y => n100);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(15), A2 => n3, B1 => 
                           data_tx_pl_15_port, B2 => n10, Y => n99);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(16), A2 => n3, B1 => 
                           data_tx_pl_16_port, B2 => n8, Y => n98);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(17), A2 => n3, B1 => 
                           data_tx_pl_17_port, B2 => n8, Y => n97);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(18), A2 => n3, B1 => 
                           data_tx_pl_18_port, B2 => n8, Y => n96);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(19), A2 => n3, B1 => 
                           data_tx_pl_19_port, B2 => n8, Y => n95);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(20), A2 => n3, B1 => 
                           data_tx_pl_20_port, B2 => n8, Y => n94);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(21), A2 => n3, B1 => 
                           data_tx_pl_21_port, B2 => n8, Y => n93);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(22), A2 => n3, B1 => 
                           data_tx_pl_22_port, B2 => n8, Y => n92);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(23), A2 => n3, B1 => 
                           data_tx_pl_23_port, B2 => n8, Y => n91);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(24), A2 => n3, B1 => 
                           data_tx_pl_24_port, B2 => n8, Y => n90);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(25), A2 => n3, B1 => 
                           data_tx_pl_25_port, B2 => n8, Y => n89);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(26), A2 => n3, B1 => 
                           data_tx_pl_26_port, B2 => n8, Y => n88);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(27), A2 => n3, B1 => 
                           data_tx_pl_27_port, B2 => n8, Y => n87);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(28), A2 => n3, B1 => 
                           data_tx_pl_28_port, B2 => n6, Y => n86);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(29), A2 => n3, B1 => 
                           data_tx_pl_29_port, B2 => n6, Y => n85);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(30), A2 => n3, B1 => 
                           data_tx_pl_30_port, B2 => n6, Y => n84);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(31), A2 => n3, B1 => 
                           data_tx_pl_31_port, B2 => n6, Y => n83);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(32), A2 => n3, B1 => 
                           data_tx_pl_32_port, B2 => n6, Y => n82);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(33), A2 => n3, B1 => 
                           data_tx_pl_33_port, B2 => n6, Y => n81);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(34), A2 => n3, B1 => 
                           data_tx_pl_34_port, B2 => n6, Y => n80);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(35), A2 => n3, B1 => 
                           data_tx_pl_35_port, B2 => n6, Y => n79);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(36), A2 => n3, B1 => 
                           data_tx_pl_36_port, B2 => n6, Y => n78);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(37), A2 => n3, B1 => 
                           data_tx_pl_37_port, B2 => n6, Y => n76);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(38), A2 => n3, B1 => 
                           data_tx_pl_38_port, B2 => n6, Y => n74);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(39), A2 => n3, B1 => 
                           data_tx_pl_39_port, B2 => n6, Y => n72);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(40), A2 => n3, B1 => 
                           data_tx_pl_40_port, B2 => n5, Y => n70);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(41), A2 => n3, B1 => 
                           data_tx_pl_41_port, B2 => n5, Y => n68);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(42), A2 => n3, B1 => 
                           data_tx_pl_42_port, B2 => n5, Y => n66);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(43), A2 => n3, B1 => 
                           data_tx_pl_43_port, B2 => n5, Y => n64);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(44), A2 => n3, B1 => 
                           data_tx_pl_44_port, B2 => n5, Y => n62);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(45), A2 => n3, B1 => 
                           data_tx_pl_45_port, B2 => n5, Y => n60);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(46), A2 => n3, B1 => 
                           data_tx_pl_46_port, B2 => n5, Y => n58);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(47), A2 => n3, B1 => 
                           data_tx_pl_47_port, B2 => n5, Y => n56);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(48), A2 => n3, B1 => 
                           data_tx_pl_48_port, B2 => n5, Y => n54);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(49), A2 => n3, B1 => 
                           data_tx_pl_49_port, B2 => n5, Y => n52);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(50), A2 => n3, B1 => 
                           data_tx_pl_50_port, B2 => n5, Y => n50);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(51), A2 => n3, B1 => 
                           data_tx_pl_51_port, B2 => n5, Y => n48);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(52), A2 => n3, B1 => 
                           data_tx_pl_52_port, B2 => n4, Y => n46);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(53), A2 => n3, B1 => 
                           data_tx_pl_53_port, B2 => n4, Y => n44);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(54), A2 => n3, B1 => 
                           data_tx_pl_54_port, B2 => n4, Y => n42);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(55), A2 => n3, B1 => 
                           data_tx_pl_55_port, B2 => n4, Y => n40);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(56), A2 => n3, B1 => 
                           data_tx_pl_56_port, B2 => n4, Y => n38);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(57), A2 => n3, B1 => 
                           data_tx_pl_57_port, B2 => n4, Y => n36);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(58), A2 => n3, B1 => 
                           data_tx_pl_58_port, B2 => n4, Y => n34);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(59), A2 => n3, B1 => 
                           data_tx_pl_59_port, B2 => n4, Y => n32);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(60), A2 => n3, B1 => 
                           data_tx_pl_60_port, B2 => n4, Y => n30);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(61), A2 => n3, B1 => 
                           data_tx_pl_61_port, B2 => n4, Y => n28);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(62), A2 => n3, B1 => 
                           data_tx_pl_62_port, B2 => n4, Y => n26);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(63), A2 => n3, B1 => 
                           data_tx_pl_63_port, B2 => n4, Y => n24);
   U68 : NAND2xp5_ASAP7_75t_R port map( A => n20, B => n22, Y => n115);
   vc_write_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n22, CLK
                           => clk, RESET => n16, SET => n1, QN => 
                           vc_write_tx_pl(0));
   vc_write_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n20, CLK
                           => clk, RESET => n16, SET => n1, QN => 
                           vc_write_tx_pl(1));
   incr_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n14, CLK => 
                           clk, RESET => n16, SET => n1, QN => incr_tx_pl(1));
   incr_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n18, CLK => 
                           clk, RESET => n16, SET => n1, QN => incr_tx_pl(0));
   data_tx_pl_reg_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n50, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_50_port);
   data_tx_pl_reg_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n52, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_49_port);
   data_tx_pl_reg_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n54, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_48_port);
   data_tx_pl_reg_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n56, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_47_port);
   data_tx_pl_reg_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n58, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_46_port);
   data_tx_pl_reg_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n60, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_45_port);
   data_tx_pl_reg_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n62, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_44_port);
   data_tx_pl_reg_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n64, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_43_port);
   data_tx_pl_reg_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n66, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_42_port);
   data_tx_pl_reg_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n68, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_41_port);
   data_tx_pl_reg_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n70, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_40_port);
   data_tx_pl_reg_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n72, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_39_port);
   data_tx_pl_reg_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n74, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_38_port);
   data_tx_pl_reg_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n76, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_37_port);
   data_tx_pl_reg_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n78, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_36_port);
   data_tx_pl_reg_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_35_port);
   data_tx_pl_reg_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n80, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_34_port);
   data_tx_pl_reg_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_33_port);
   data_tx_pl_reg_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n82, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_32_port);
   data_tx_pl_reg_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_31_port);
   data_tx_pl_reg_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n84, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_30_port);
   data_tx_pl_reg_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n102, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_12_port);
   data_tx_pl_reg_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_11_port);
   data_tx_pl_reg_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n104, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_10_port);
   data_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n114, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_0_port);
   data_tx_pl_reg_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n24, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_63_port);
   data_tx_pl_reg_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n26, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_62_port);
   data_tx_pl_reg_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n28, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_61_port);
   data_tx_pl_reg_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n30, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_60_port);
   data_tx_pl_reg_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n32, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_59_port);
   data_tx_pl_reg_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n34, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_58_port);
   data_tx_pl_reg_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n36, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_57_port);
   data_tx_pl_reg_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n38, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_56_port);
   data_tx_pl_reg_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n40, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_55_port);
   data_tx_pl_reg_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n42, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_54_port);
   data_tx_pl_reg_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n44, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_53_port);
   data_tx_pl_reg_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n46, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_52_port);
   data_tx_pl_reg_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n48, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_51_port);
   data_tx_pl_reg_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_29_port);
   data_tx_pl_reg_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n86, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_28_port);
   data_tx_pl_reg_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_27_port);
   data_tx_pl_reg_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n88, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_26_port);
   data_tx_pl_reg_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_25_port);
   data_tx_pl_reg_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n90, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_24_port);
   data_tx_pl_reg_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_23_port);
   data_tx_pl_reg_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n92, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_22_port);
   data_tx_pl_reg_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_21_port);
   data_tx_pl_reg_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n94, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_20_port);
   data_tx_pl_reg_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_19_port);
   data_tx_pl_reg_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n96, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_18_port);
   data_tx_pl_reg_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_17_port);
   data_tx_pl_reg_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n98, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_16_port);
   data_tx_pl_reg_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_15_port);
   data_tx_pl_reg_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n100, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_14_port);
   data_tx_pl_reg_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_13_port);
   data_tx_pl_reg_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_9_port);
   data_tx_pl_reg_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n106, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_8_port);
   data_tx_pl_reg_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_7_port);
   data_tx_pl_reg_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n108, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_6_port);
   data_tx_pl_reg_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_5_port);
   data_tx_pl_reg_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n110, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_4_port);
   data_tx_pl_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_3_port);
   data_tx_pl_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n112, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_2_port);
   data_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_1_port);
   U67 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U69 : INVx2_ASAP7_75t_R port map( A => rst, Y => n16);
   U70 : INVx1_ASAP7_75t_R port map( A => n12, Y => n3);
   U71 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n12);
   U72 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n10);
   U73 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n8);
   U74 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n6);
   U75 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n5);
   U76 : HB1xp67_ASAP7_75t_R port map( A => n115, Y => n4);
   U77 : INVx1_ASAP7_75t_R port map( A => incr_tx(1), Y => n14);
   U78 : INVx1_ASAP7_75t_R port map( A => incr_tx(0), Y => n18);
   U79 : INVx1_ASAP7_75t_R port map( A => vc_write_tx(1), Y => n20);
   U80 : INVx1_ASAP7_75t_R port map( A => vc_write_tx(0), Y => n22);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity vc_input_buffer_2_0000000200000002_5 is

   port( clk, rst : in std_logic;  data_rx : in std_logic_vector (63 downto 0);
         vc_write_rx, vc_transfer : in std_logic_vector (1 downto 0);  
         valid_data_vc : out std_logic_vector (1 downto 0);  data_transfer : 
         out std_logic_vector (63 downto 0);  header : out std_logic_vector (19
         downto 0));

end vc_input_buffer_2_0000000200000002_5;

architecture SYN_rtl of vc_input_buffer_2_0000000200000002_5 is

   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component fifo_buff_depth2_9
      port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, 
            clk, rst : in std_logic;  data_out : out std_logic_vector (63 
            downto 0);  valid_data : out std_logic);
   end component;
   
   component fifo_buff_depth2_10
      port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, 
            clk, rst : in std_logic;  data_out : out std_logic_vector (63 
            downto 0);  valid_data : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal header_1_PACKET_LENGTH_3_port, header_1_PACKET_LENGTH_2_port, 
      header_1_PACKET_LENGTH_1_port, header_1_PACKET_LENGTH_0_port, 
      header_1_X_DEST_1_port, header_1_X_DEST_0_port, header_1_Y_DEST_1_port, 
      header_1_Y_DEST_0_port, header_1_Z_DEST_1_port, header_1_Z_DEST_0_port, 
      header_0_PACKET_LENGTH_3_port, header_0_PACKET_LENGTH_2_port, 
      header_0_PACKET_LENGTH_1_port, header_0_PACKET_LENGTH_0_port, 
      header_0_X_DEST_1_port, header_0_X_DEST_0_port, header_0_Y_DEST_1_port, 
      header_0_Y_DEST_0_port, header_0_Z_DEST_1_port, header_0_Z_DEST_0_port, 
      buffer_out_vector_1_63_port, buffer_out_vector_1_62_port, 
      buffer_out_vector_1_61_port, buffer_out_vector_1_60_port, 
      buffer_out_vector_1_59_port, buffer_out_vector_1_58_port, 
      buffer_out_vector_1_57_port, buffer_out_vector_1_56_port, 
      buffer_out_vector_1_55_port, buffer_out_vector_1_54_port, 
      buffer_out_vector_1_53_port, buffer_out_vector_1_52_port, 
      buffer_out_vector_1_51_port, buffer_out_vector_1_50_port, 
      buffer_out_vector_1_49_port, buffer_out_vector_1_48_port, 
      buffer_out_vector_1_47_port, buffer_out_vector_1_46_port, 
      buffer_out_vector_1_45_port, buffer_out_vector_1_44_port, 
      buffer_out_vector_1_43_port, buffer_out_vector_1_42_port, 
      buffer_out_vector_1_41_port, buffer_out_vector_1_40_port, 
      buffer_out_vector_1_39_port, buffer_out_vector_1_38_port, 
      buffer_out_vector_1_37_port, buffer_out_vector_1_36_port, 
      buffer_out_vector_1_35_port, buffer_out_vector_1_34_port, 
      buffer_out_vector_1_33_port, buffer_out_vector_1_32_port, 
      buffer_out_vector_1_31_port, buffer_out_vector_1_30_port, 
      buffer_out_vector_1_29_port, buffer_out_vector_1_28_port, 
      buffer_out_vector_1_27_port, buffer_out_vector_1_26_port, 
      buffer_out_vector_1_25_port, buffer_out_vector_1_24_port, 
      buffer_out_vector_1_23_port, buffer_out_vector_1_22_port, 
      buffer_out_vector_1_21_port, buffer_out_vector_1_20_port, 
      buffer_out_vector_1_19_port, buffer_out_vector_1_18_port, 
      buffer_out_vector_1_17_port, buffer_out_vector_1_16_port, 
      buffer_out_vector_1_15_port, buffer_out_vector_1_14_port, 
      buffer_out_vector_1_13_port, buffer_out_vector_1_12_port, 
      buffer_out_vector_1_11_port, buffer_out_vector_1_10_port, 
      buffer_out_vector_0_63_port, buffer_out_vector_0_62_port, 
      buffer_out_vector_0_61_port, buffer_out_vector_0_60_port, 
      buffer_out_vector_0_59_port, buffer_out_vector_0_58_port, 
      buffer_out_vector_0_57_port, buffer_out_vector_0_56_port, 
      buffer_out_vector_0_55_port, buffer_out_vector_0_54_port, 
      buffer_out_vector_0_53_port, buffer_out_vector_0_52_port, 
      buffer_out_vector_0_51_port, buffer_out_vector_0_50_port, 
      buffer_out_vector_0_49_port, buffer_out_vector_0_48_port, 
      buffer_out_vector_0_47_port, buffer_out_vector_0_46_port, 
      buffer_out_vector_0_45_port, buffer_out_vector_0_44_port, 
      buffer_out_vector_0_43_port, buffer_out_vector_0_42_port, 
      buffer_out_vector_0_41_port, buffer_out_vector_0_40_port, 
      buffer_out_vector_0_39_port, buffer_out_vector_0_38_port, 
      buffer_out_vector_0_37_port, buffer_out_vector_0_36_port, 
      buffer_out_vector_0_35_port, buffer_out_vector_0_34_port, 
      buffer_out_vector_0_33_port, buffer_out_vector_0_32_port, 
      buffer_out_vector_0_31_port, buffer_out_vector_0_30_port, 
      buffer_out_vector_0_29_port, buffer_out_vector_0_28_port, 
      buffer_out_vector_0_27_port, buffer_out_vector_0_26_port, 
      buffer_out_vector_0_25_port, buffer_out_vector_0_24_port, 
      buffer_out_vector_0_23_port, buffer_out_vector_0_22_port, 
      buffer_out_vector_0_21_port, buffer_out_vector_0_20_port, 
      buffer_out_vector_0_19_port, buffer_out_vector_0_18_port, 
      buffer_out_vector_0_17_port, buffer_out_vector_0_16_port, 
      buffer_out_vector_0_15_port, buffer_out_vector_0_14_port, 
      buffer_out_vector_0_13_port, buffer_out_vector_0_12_port, 
      buffer_out_vector_0_11_port, buffer_out_vector_0_10_port, n1, n2, n3, n4,
      n5, n6, n7, n8 : std_logic;

begin
   header <= ( header_1_PACKET_LENGTH_3_port, header_1_PACKET_LENGTH_2_port, 
      header_1_PACKET_LENGTH_1_port, header_1_PACKET_LENGTH_0_port, 
      header_1_X_DEST_1_port, header_1_X_DEST_0_port, header_1_Y_DEST_1_port, 
      header_1_Y_DEST_0_port, header_1_Z_DEST_1_port, header_1_Z_DEST_0_port, 
      header_0_PACKET_LENGTH_3_port, header_0_PACKET_LENGTH_2_port, 
      header_0_PACKET_LENGTH_1_port, header_0_PACKET_LENGTH_0_port, 
      header_0_X_DEST_1_port, header_0_X_DEST_0_port, header_0_Y_DEST_1_port, 
      header_0_Y_DEST_0_port, header_0_Z_DEST_1_port, header_0_Z_DEST_0_port );
   
   U2 : AO22x1_ASAP7_75t_R port map( A1 => n3, A2 => 
                           buffer_out_vector_1_30_port, B1 => 
                           buffer_out_vector_0_30_port, B2 => n4, Y => 
                           data_transfer(30));
   U3 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_31_port, A2 => 
                           n3, B1 => buffer_out_vector_0_31_port, B2 => n4, Y 
                           => data_transfer(31));
   U4 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_32_port, A2 => 
                           n3, B1 => buffer_out_vector_0_32_port, B2 => n4, Y 
                           => data_transfer(32));
   U5 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_33_port, A2 => 
                           n3, B1 => buffer_out_vector_0_33_port, B2 => n4, Y 
                           => data_transfer(33));
   U6 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_34_port, A2 => 
                           n3, B1 => buffer_out_vector_0_34_port, B2 => n4, Y 
                           => data_transfer(34));
   U7 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_35_port, A2 => 
                           n3, B1 => buffer_out_vector_0_35_port, B2 => n6, Y 
                           => data_transfer(35));
   U8 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_36_port, A2 => 
                           n3, B1 => buffer_out_vector_0_36_port, B2 => n5, Y 
                           => data_transfer(36));
   U9 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_37_port, A2 => 
                           n3, B1 => buffer_out_vector_0_37_port, B2 => n7, Y 
                           => data_transfer(37));
   U10 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_38_port, A2 => 
                           n3, B1 => buffer_out_vector_0_38_port, B2 => n6, Y 
                           => data_transfer(38));
   U11 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_39_port, A2 => 
                           n3, B1 => buffer_out_vector_0_39_port, B2 => n5, Y 
                           => data_transfer(39));
   U12 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_40_port, A2 => 
                           n3, B1 => buffer_out_vector_0_40_port, B2 => n7, Y 
                           => data_transfer(40));
   U13 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_41_port, A2 => 
                           n3, B1 => buffer_out_vector_0_41_port, B2 => n6, Y 
                           => data_transfer(41));
   U14 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_42_port, A2 => 
                           n3, B1 => buffer_out_vector_0_42_port, B2 => n5, Y 
                           => data_transfer(42));
   U15 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_43_port, A2 => 
                           n3, B1 => buffer_out_vector_0_43_port, B2 => n7, Y 
                           => data_transfer(43));
   U16 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_44_port, A2 => 
                           n3, B1 => buffer_out_vector_0_44_port, B2 => n7, Y 
                           => data_transfer(44));
   U17 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_45_port, A2 => 
                           n3, B1 => buffer_out_vector_0_45_port, B2 => n6, Y 
                           => data_transfer(45));
   U18 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_46_port, A2 => 
                           n3, B1 => buffer_out_vector_0_46_port, B2 => n5, Y 
                           => data_transfer(46));
   U19 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_47_port, A2 => 
                           n3, B1 => buffer_out_vector_0_47_port, B2 => n6, Y 
                           => data_transfer(47));
   U20 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_48_port, A2 => 
                           n3, B1 => buffer_out_vector_0_48_port, B2 => n6, Y 
                           => data_transfer(48));
   U21 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_49_port, A2 => 
                           n3, B1 => buffer_out_vector_0_49_port, B2 => n7, Y 
                           => data_transfer(49));
   U22 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_50_port, A2 => 
                           n3, B1 => buffer_out_vector_0_50_port, B2 => n6, Y 
                           => data_transfer(50));
   U23 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_51_port, A2 => 
                           n2, B1 => buffer_out_vector_0_51_port, B2 => n7, Y 
                           => data_transfer(51));
   U24 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_52_port, A2 => 
                           n2, B1 => buffer_out_vector_0_52_port, B2 => n5, Y 
                           => data_transfer(52));
   U25 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_53_port, A2 => 
                           n2, B1 => buffer_out_vector_0_53_port, B2 => n6, Y 
                           => data_transfer(53));
   U26 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_54_port, A2 => 
                           n2, B1 => buffer_out_vector_0_54_port, B2 => n7, Y 
                           => data_transfer(54));
   U27 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_55_port, A2 => 
                           n2, B1 => buffer_out_vector_0_55_port, B2 => n6, Y 
                           => data_transfer(55));
   U28 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_56_port, A2 => 
                           n2, B1 => buffer_out_vector_0_56_port, B2 => n5, Y 
                           => data_transfer(56));
   U29 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_57_port, A2 => 
                           n2, B1 => buffer_out_vector_0_57_port, B2 => n7, Y 
                           => data_transfer(57));
   U30 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_58_port, A2 => 
                           n2, B1 => buffer_out_vector_0_58_port, B2 => n6, Y 
                           => data_transfer(58));
   U31 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_59_port, A2 => 
                           n2, B1 => buffer_out_vector_0_59_port, B2 => n5, Y 
                           => data_transfer(59));
   U32 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_60_port, A2 => 
                           n2, B1 => buffer_out_vector_0_60_port, B2 => n6, Y 
                           => data_transfer(60));
   U33 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_61_port, A2 => 
                           n2, B1 => buffer_out_vector_0_61_port, B2 => n7, Y 
                           => data_transfer(61));
   U34 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_62_port, A2 => 
                           n2, B1 => buffer_out_vector_0_62_port, B2 => n6, Y 
                           => data_transfer(62));
   U35 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_63_port, A2 => 
                           n2, B1 => buffer_out_vector_0_63_port, B2 => n5, Y 
                           => data_transfer(63));
   U36 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_0_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_0_port, B2 => n7
                           , Y => data_transfer(0));
   U37 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_1_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_1_port, B2 => n5
                           , Y => data_transfer(1));
   U38 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_2_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_2_port, B2 => n7
                           , Y => data_transfer(2));
   U39 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_3_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_3_port, B2 => n5
                           , Y => data_transfer(3));
   U40 : AO22x1_ASAP7_75t_R port map( A1 => header_1_X_DEST_0_port, A2 => n2, 
                           B1 => header_0_X_DEST_0_port, B2 => n5, Y => 
                           data_transfer(4));
   U41 : AO22x1_ASAP7_75t_R port map( A1 => header_1_X_DEST_1_port, A2 => n2, 
                           B1 => header_0_X_DEST_1_port, B2 => n5, Y => 
                           data_transfer(5));
   U42 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Y_DEST_0_port, A2 => n2, 
                           B1 => header_0_Y_DEST_0_port, B2 => n5, Y => 
                           data_transfer(6));
   U43 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Y_DEST_1_port, A2 => n2, 
                           B1 => header_0_Y_DEST_1_port, B2 => n5, Y => 
                           data_transfer(7));
   U44 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Z_DEST_0_port, A2 => n2, 
                           B1 => header_0_Z_DEST_0_port, B2 => n5, Y => 
                           data_transfer(8));
   U45 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Z_DEST_1_port, A2 => n2, 
                           B1 => header_0_Z_DEST_1_port, B2 => n5, Y => 
                           data_transfer(9));
   U46 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_10_port, A2 => 
                           n2, B1 => buffer_out_vector_0_10_port, B2 => n5, Y 
                           => data_transfer(10));
   U47 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_11_port, A2 => 
                           n2, B1 => buffer_out_vector_0_11_port, B2 => n6, Y 
                           => data_transfer(11));
   U48 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_12_port, A2 => 
                           n2, B1 => buffer_out_vector_0_12_port, B2 => n6, Y 
                           => data_transfer(12));
   U49 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_13_port, A2 => 
                           n2, B1 => buffer_out_vector_0_13_port, B2 => n6, Y 
                           => data_transfer(13));
   U50 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_14_port, A2 => 
                           n2, B1 => buffer_out_vector_0_14_port, B2 => n6, Y 
                           => data_transfer(14));
   U51 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_15_port, A2 => 
                           n2, B1 => buffer_out_vector_0_15_port, B2 => n6, Y 
                           => data_transfer(15));
   U52 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_16_port, A2 => 
                           n2, B1 => buffer_out_vector_0_16_port, B2 => n6, Y 
                           => data_transfer(16));
   U53 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_17_port, A2 => 
                           n2, B1 => buffer_out_vector_0_17_port, B2 => n6, Y 
                           => data_transfer(17));
   U54 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_18_port, A2 => 
                           n2, B1 => buffer_out_vector_0_18_port, B2 => n6, Y 
                           => data_transfer(18));
   U55 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_19_port, A2 => 
                           n2, B1 => buffer_out_vector_0_19_port, B2 => n7, Y 
                           => data_transfer(19));
   U56 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_20_port, A2 => 
                           n2, B1 => buffer_out_vector_0_20_port, B2 => n7, Y 
                           => data_transfer(20));
   U57 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_21_port, A2 => 
                           n2, B1 => buffer_out_vector_0_21_port, B2 => n7, Y 
                           => data_transfer(21));
   U58 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_22_port, A2 => 
                           n2, B1 => buffer_out_vector_0_22_port, B2 => n7, Y 
                           => data_transfer(22));
   U59 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_23_port, A2 => 
                           n2, B1 => buffer_out_vector_0_23_port, B2 => n7, Y 
                           => data_transfer(23));
   U60 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_24_port, A2 => 
                           n2, B1 => buffer_out_vector_0_24_port, B2 => n7, Y 
                           => data_transfer(24));
   U61 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_25_port, A2 => 
                           n2, B1 => buffer_out_vector_0_25_port, B2 => n7, Y 
                           => data_transfer(25));
   U62 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_26_port, A2 => 
                           n2, B1 => buffer_out_vector_0_26_port, B2 => n7, Y 
                           => data_transfer(26));
   U63 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_27_port, A2 => 
                           n2, B1 => buffer_out_vector_0_27_port, B2 => n5, Y 
                           => data_transfer(27));
   U64 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_28_port, A2 => 
                           n2, B1 => buffer_out_vector_0_28_port, B2 => n5, Y 
                           => data_transfer(28));
   U65 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_29_port, A2 => 
                           n2, B1 => buffer_out_vector_0_29_port, B2 => n5, Y 
                           => data_transfer(29));
   fifo_i_0 : fifo_buff_depth2_10 port map( data_in(63) => data_rx(63), 
                           data_in(62) => data_rx(62), data_in(61) => 
                           data_rx(61), data_in(60) => data_rx(60), data_in(59)
                           => data_rx(59), data_in(58) => data_rx(58), 
                           data_in(57) => data_rx(57), data_in(56) => 
                           data_rx(56), data_in(55) => data_rx(55), data_in(54)
                           => data_rx(54), data_in(53) => data_rx(53), 
                           data_in(52) => data_rx(52), data_in(51) => 
                           data_rx(51), data_in(50) => data_rx(50), data_in(49)
                           => data_rx(49), data_in(48) => data_rx(48), 
                           data_in(47) => data_rx(47), data_in(46) => 
                           data_rx(46), data_in(45) => data_rx(45), data_in(44)
                           => data_rx(44), data_in(43) => data_rx(43), 
                           data_in(42) => data_rx(42), data_in(41) => 
                           data_rx(41), data_in(40) => data_rx(40), data_in(39)
                           => data_rx(39), data_in(38) => data_rx(38), 
                           data_in(37) => data_rx(37), data_in(36) => 
                           data_rx(36), data_in(35) => data_rx(35), data_in(34)
                           => data_rx(34), data_in(33) => data_rx(33), 
                           data_in(32) => data_rx(32), data_in(31) => 
                           data_rx(31), data_in(30) => data_rx(30), data_in(29)
                           => data_rx(29), data_in(28) => data_rx(28), 
                           data_in(27) => data_rx(27), data_in(26) => 
                           data_rx(26), data_in(25) => data_rx(25), data_in(24)
                           => data_rx(24), data_in(23) => data_rx(23), 
                           data_in(22) => data_rx(22), data_in(21) => 
                           data_rx(21), data_in(20) => data_rx(20), data_in(19)
                           => data_rx(19), data_in(18) => data_rx(18), 
                           data_in(17) => data_rx(17), data_in(16) => 
                           data_rx(16), data_in(15) => data_rx(15), data_in(14)
                           => data_rx(14), data_in(13) => data_rx(13), 
                           data_in(12) => data_rx(12), data_in(11) => 
                           data_rx(11), data_in(10) => data_rx(10), data_in(9) 
                           => data_rx(9), data_in(8) => data_rx(8), data_in(7) 
                           => data_rx(7), data_in(6) => data_rx(6), data_in(5) 
                           => data_rx(5), data_in(4) => data_rx(4), data_in(3) 
                           => data_rx(3), data_in(2) => data_rx(2), data_in(1) 
                           => data_rx(1), data_in(0) => data_rx(0), write_en =>
                           vc_write_rx(0), read_en => vc_transfer(0), clk => 
                           clk, rst => n8, data_out(63) => 
                           buffer_out_vector_0_63_port, data_out(62) => 
                           buffer_out_vector_0_62_port, data_out(61) => 
                           buffer_out_vector_0_61_port, data_out(60) => 
                           buffer_out_vector_0_60_port, data_out(59) => 
                           buffer_out_vector_0_59_port, data_out(58) => 
                           buffer_out_vector_0_58_port, data_out(57) => 
                           buffer_out_vector_0_57_port, data_out(56) => 
                           buffer_out_vector_0_56_port, data_out(55) => 
                           buffer_out_vector_0_55_port, data_out(54) => 
                           buffer_out_vector_0_54_port, data_out(53) => 
                           buffer_out_vector_0_53_port, data_out(52) => 
                           buffer_out_vector_0_52_port, data_out(51) => 
                           buffer_out_vector_0_51_port, data_out(50) => 
                           buffer_out_vector_0_50_port, data_out(49) => 
                           buffer_out_vector_0_49_port, data_out(48) => 
                           buffer_out_vector_0_48_port, data_out(47) => 
                           buffer_out_vector_0_47_port, data_out(46) => 
                           buffer_out_vector_0_46_port, data_out(45) => 
                           buffer_out_vector_0_45_port, data_out(44) => 
                           buffer_out_vector_0_44_port, data_out(43) => 
                           buffer_out_vector_0_43_port, data_out(42) => 
                           buffer_out_vector_0_42_port, data_out(41) => 
                           buffer_out_vector_0_41_port, data_out(40) => 
                           buffer_out_vector_0_40_port, data_out(39) => 
                           buffer_out_vector_0_39_port, data_out(38) => 
                           buffer_out_vector_0_38_port, data_out(37) => 
                           buffer_out_vector_0_37_port, data_out(36) => 
                           buffer_out_vector_0_36_port, data_out(35) => 
                           buffer_out_vector_0_35_port, data_out(34) => 
                           buffer_out_vector_0_34_port, data_out(33) => 
                           buffer_out_vector_0_33_port, data_out(32) => 
                           buffer_out_vector_0_32_port, data_out(31) => 
                           buffer_out_vector_0_31_port, data_out(30) => 
                           buffer_out_vector_0_30_port, data_out(29) => 
                           buffer_out_vector_0_29_port, data_out(28) => 
                           buffer_out_vector_0_28_port, data_out(27) => 
                           buffer_out_vector_0_27_port, data_out(26) => 
                           buffer_out_vector_0_26_port, data_out(25) => 
                           buffer_out_vector_0_25_port, data_out(24) => 
                           buffer_out_vector_0_24_port, data_out(23) => 
                           buffer_out_vector_0_23_port, data_out(22) => 
                           buffer_out_vector_0_22_port, data_out(21) => 
                           buffer_out_vector_0_21_port, data_out(20) => 
                           buffer_out_vector_0_20_port, data_out(19) => 
                           buffer_out_vector_0_19_port, data_out(18) => 
                           buffer_out_vector_0_18_port, data_out(17) => 
                           buffer_out_vector_0_17_port, data_out(16) => 
                           buffer_out_vector_0_16_port, data_out(15) => 
                           buffer_out_vector_0_15_port, data_out(14) => 
                           buffer_out_vector_0_14_port, data_out(13) => 
                           buffer_out_vector_0_13_port, data_out(12) => 
                           buffer_out_vector_0_12_port, data_out(11) => 
                           buffer_out_vector_0_11_port, data_out(10) => 
                           buffer_out_vector_0_10_port, data_out(9) => 
                           header_0_Z_DEST_1_port, data_out(8) => 
                           header_0_Z_DEST_0_port, data_out(7) => 
                           header_0_Y_DEST_1_port, data_out(6) => 
                           header_0_Y_DEST_0_port, data_out(5) => 
                           header_0_X_DEST_1_port, data_out(4) => 
                           header_0_X_DEST_0_port, data_out(3) => 
                           header_0_PACKET_LENGTH_3_port, data_out(2) => 
                           header_0_PACKET_LENGTH_2_port, data_out(1) => 
                           header_0_PACKET_LENGTH_1_port, data_out(0) => 
                           header_0_PACKET_LENGTH_0_port, valid_data => 
                           valid_data_vc(0));
   fifo_i_1 : fifo_buff_depth2_9 port map( data_in(63) => data_rx(63), 
                           data_in(62) => data_rx(62), data_in(61) => 
                           data_rx(61), data_in(60) => data_rx(60), data_in(59)
                           => data_rx(59), data_in(58) => data_rx(58), 
                           data_in(57) => data_rx(57), data_in(56) => 
                           data_rx(56), data_in(55) => data_rx(55), data_in(54)
                           => data_rx(54), data_in(53) => data_rx(53), 
                           data_in(52) => data_rx(52), data_in(51) => 
                           data_rx(51), data_in(50) => data_rx(50), data_in(49)
                           => data_rx(49), data_in(48) => data_rx(48), 
                           data_in(47) => data_rx(47), data_in(46) => 
                           data_rx(46), data_in(45) => data_rx(45), data_in(44)
                           => data_rx(44), data_in(43) => data_rx(43), 
                           data_in(42) => data_rx(42), data_in(41) => 
                           data_rx(41), data_in(40) => data_rx(40), data_in(39)
                           => data_rx(39), data_in(38) => data_rx(38), 
                           data_in(37) => data_rx(37), data_in(36) => 
                           data_rx(36), data_in(35) => data_rx(35), data_in(34)
                           => data_rx(34), data_in(33) => data_rx(33), 
                           data_in(32) => data_rx(32), data_in(31) => 
                           data_rx(31), data_in(30) => data_rx(30), data_in(29)
                           => data_rx(29), data_in(28) => data_rx(28), 
                           data_in(27) => data_rx(27), data_in(26) => 
                           data_rx(26), data_in(25) => data_rx(25), data_in(24)
                           => data_rx(24), data_in(23) => data_rx(23), 
                           data_in(22) => data_rx(22), data_in(21) => 
                           data_rx(21), data_in(20) => data_rx(20), data_in(19)
                           => data_rx(19), data_in(18) => data_rx(18), 
                           data_in(17) => data_rx(17), data_in(16) => 
                           data_rx(16), data_in(15) => data_rx(15), data_in(14)
                           => data_rx(14), data_in(13) => data_rx(13), 
                           data_in(12) => data_rx(12), data_in(11) => 
                           data_rx(11), data_in(10) => data_rx(10), data_in(9) 
                           => data_rx(9), data_in(8) => data_rx(8), data_in(7) 
                           => data_rx(7), data_in(6) => data_rx(6), data_in(5) 
                           => data_rx(5), data_in(4) => data_rx(4), data_in(3) 
                           => data_rx(3), data_in(2) => data_rx(2), data_in(1) 
                           => data_rx(1), data_in(0) => data_rx(0), write_en =>
                           vc_write_rx(1), read_en => n2, clk => clk, rst => n8
                           , data_out(63) => buffer_out_vector_1_63_port, 
                           data_out(62) => buffer_out_vector_1_62_port, 
                           data_out(61) => buffer_out_vector_1_61_port, 
                           data_out(60) => buffer_out_vector_1_60_port, 
                           data_out(59) => buffer_out_vector_1_59_port, 
                           data_out(58) => buffer_out_vector_1_58_port, 
                           data_out(57) => buffer_out_vector_1_57_port, 
                           data_out(56) => buffer_out_vector_1_56_port, 
                           data_out(55) => buffer_out_vector_1_55_port, 
                           data_out(54) => buffer_out_vector_1_54_port, 
                           data_out(53) => buffer_out_vector_1_53_port, 
                           data_out(52) => buffer_out_vector_1_52_port, 
                           data_out(51) => buffer_out_vector_1_51_port, 
                           data_out(50) => buffer_out_vector_1_50_port, 
                           data_out(49) => buffer_out_vector_1_49_port, 
                           data_out(48) => buffer_out_vector_1_48_port, 
                           data_out(47) => buffer_out_vector_1_47_port, 
                           data_out(46) => buffer_out_vector_1_46_port, 
                           data_out(45) => buffer_out_vector_1_45_port, 
                           data_out(44) => buffer_out_vector_1_44_port, 
                           data_out(43) => buffer_out_vector_1_43_port, 
                           data_out(42) => buffer_out_vector_1_42_port, 
                           data_out(41) => buffer_out_vector_1_41_port, 
                           data_out(40) => buffer_out_vector_1_40_port, 
                           data_out(39) => buffer_out_vector_1_39_port, 
                           data_out(38) => buffer_out_vector_1_38_port, 
                           data_out(37) => buffer_out_vector_1_37_port, 
                           data_out(36) => buffer_out_vector_1_36_port, 
                           data_out(35) => buffer_out_vector_1_35_port, 
                           data_out(34) => buffer_out_vector_1_34_port, 
                           data_out(33) => buffer_out_vector_1_33_port, 
                           data_out(32) => buffer_out_vector_1_32_port, 
                           data_out(31) => buffer_out_vector_1_31_port, 
                           data_out(30) => buffer_out_vector_1_30_port, 
                           data_out(29) => buffer_out_vector_1_29_port, 
                           data_out(28) => buffer_out_vector_1_28_port, 
                           data_out(27) => buffer_out_vector_1_27_port, 
                           data_out(26) => buffer_out_vector_1_26_port, 
                           data_out(25) => buffer_out_vector_1_25_port, 
                           data_out(24) => buffer_out_vector_1_24_port, 
                           data_out(23) => buffer_out_vector_1_23_port, 
                           data_out(22) => buffer_out_vector_1_22_port, 
                           data_out(21) => buffer_out_vector_1_21_port, 
                           data_out(20) => buffer_out_vector_1_20_port, 
                           data_out(19) => buffer_out_vector_1_19_port, 
                           data_out(18) => buffer_out_vector_1_18_port, 
                           data_out(17) => buffer_out_vector_1_17_port, 
                           data_out(16) => buffer_out_vector_1_16_port, 
                           data_out(15) => buffer_out_vector_1_15_port, 
                           data_out(14) => buffer_out_vector_1_14_port, 
                           data_out(13) => buffer_out_vector_1_13_port, 
                           data_out(12) => buffer_out_vector_1_12_port, 
                           data_out(11) => buffer_out_vector_1_11_port, 
                           data_out(10) => buffer_out_vector_1_10_port, 
                           data_out(9) => header_1_Z_DEST_1_port, data_out(8) 
                           => header_1_Z_DEST_0_port, data_out(7) => 
                           header_1_Y_DEST_1_port, data_out(6) => 
                           header_1_Y_DEST_0_port, data_out(5) => 
                           header_1_X_DEST_1_port, data_out(4) => 
                           header_1_X_DEST_0_port, data_out(3) => 
                           header_1_PACKET_LENGTH_3_port, data_out(2) => 
                           header_1_PACKET_LENGTH_2_port, data_out(1) => 
                           header_1_PACKET_LENGTH_1_port, data_out(0) => 
                           header_1_PACKET_LENGTH_0_port, valid_data => 
                           valid_data_vc(1));
   U1 : INVx1_ASAP7_75t_R port map( A => n4, Y => n2);
   U66 : INVx1_ASAP7_75t_R port map( A => n4, Y => n3);
   U67 : INVx1_ASAP7_75t_R port map( A => n1, Y => n4);
   U68 : INVx1_ASAP7_75t_R port map( A => n1, Y => n5);
   U69 : INVx1_ASAP7_75t_R port map( A => n1, Y => n6);
   U70 : INVx1_ASAP7_75t_R port map( A => n1, Y => n7);
   U71 : HB1xp67_ASAP7_75t_R port map( A => vc_transfer(1), Y => n1);
   U72 : HB1xp67_ASAP7_75t_R port map( A => rst, Y => n8);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity vc_input_buffer_2_0000000200000002_4 is

   port( clk, rst : in std_logic;  data_rx : in std_logic_vector (63 downto 0);
         vc_write_rx, vc_transfer : in std_logic_vector (1 downto 0);  
         valid_data_vc : out std_logic_vector (1 downto 0);  data_transfer : 
         out std_logic_vector (63 downto 0);  header : out std_logic_vector (19
         downto 0));

end vc_input_buffer_2_0000000200000002_4;

architecture SYN_rtl of vc_input_buffer_2_0000000200000002_4 is

   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component fifo_buff_depth2_7
      port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, 
            clk, rst : in std_logic;  data_out : out std_logic_vector (63 
            downto 0);  valid_data : out std_logic);
   end component;
   
   component fifo_buff_depth2_8
      port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, 
            clk, rst : in std_logic;  data_out : out std_logic_vector (63 
            downto 0);  valid_data : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal header_1_PACKET_LENGTH_3_port, header_1_PACKET_LENGTH_2_port, 
      header_1_PACKET_LENGTH_1_port, header_1_PACKET_LENGTH_0_port, 
      header_1_X_DEST_1_port, header_1_X_DEST_0_port, header_1_Y_DEST_1_port, 
      header_1_Y_DEST_0_port, header_1_Z_DEST_1_port, header_1_Z_DEST_0_port, 
      header_0_PACKET_LENGTH_3_port, header_0_PACKET_LENGTH_2_port, 
      header_0_PACKET_LENGTH_1_port, header_0_PACKET_LENGTH_0_port, 
      header_0_X_DEST_1_port, header_0_X_DEST_0_port, header_0_Y_DEST_1_port, 
      header_0_Y_DEST_0_port, header_0_Z_DEST_1_port, header_0_Z_DEST_0_port, 
      buffer_out_vector_1_63_port, buffer_out_vector_1_62_port, 
      buffer_out_vector_1_61_port, buffer_out_vector_1_60_port, 
      buffer_out_vector_1_59_port, buffer_out_vector_1_58_port, 
      buffer_out_vector_1_57_port, buffer_out_vector_1_56_port, 
      buffer_out_vector_1_55_port, buffer_out_vector_1_54_port, 
      buffer_out_vector_1_53_port, buffer_out_vector_1_52_port, 
      buffer_out_vector_1_51_port, buffer_out_vector_1_50_port, 
      buffer_out_vector_1_49_port, buffer_out_vector_1_48_port, 
      buffer_out_vector_1_47_port, buffer_out_vector_1_46_port, 
      buffer_out_vector_1_45_port, buffer_out_vector_1_44_port, 
      buffer_out_vector_1_43_port, buffer_out_vector_1_42_port, 
      buffer_out_vector_1_41_port, buffer_out_vector_1_40_port, 
      buffer_out_vector_1_39_port, buffer_out_vector_1_38_port, 
      buffer_out_vector_1_37_port, buffer_out_vector_1_36_port, 
      buffer_out_vector_1_35_port, buffer_out_vector_1_34_port, 
      buffer_out_vector_1_33_port, buffer_out_vector_1_32_port, 
      buffer_out_vector_1_31_port, buffer_out_vector_1_30_port, 
      buffer_out_vector_1_29_port, buffer_out_vector_1_28_port, 
      buffer_out_vector_1_27_port, buffer_out_vector_1_26_port, 
      buffer_out_vector_1_25_port, buffer_out_vector_1_24_port, 
      buffer_out_vector_1_23_port, buffer_out_vector_1_22_port, 
      buffer_out_vector_1_21_port, buffer_out_vector_1_20_port, 
      buffer_out_vector_1_19_port, buffer_out_vector_1_18_port, 
      buffer_out_vector_1_17_port, buffer_out_vector_1_16_port, 
      buffer_out_vector_1_15_port, buffer_out_vector_1_14_port, 
      buffer_out_vector_1_13_port, buffer_out_vector_1_12_port, 
      buffer_out_vector_1_11_port, buffer_out_vector_1_10_port, 
      buffer_out_vector_0_63_port, buffer_out_vector_0_62_port, 
      buffer_out_vector_0_61_port, buffer_out_vector_0_60_port, 
      buffer_out_vector_0_59_port, buffer_out_vector_0_58_port, 
      buffer_out_vector_0_57_port, buffer_out_vector_0_56_port, 
      buffer_out_vector_0_55_port, buffer_out_vector_0_54_port, 
      buffer_out_vector_0_53_port, buffer_out_vector_0_52_port, 
      buffer_out_vector_0_51_port, buffer_out_vector_0_50_port, 
      buffer_out_vector_0_49_port, buffer_out_vector_0_48_port, 
      buffer_out_vector_0_47_port, buffer_out_vector_0_46_port, 
      buffer_out_vector_0_45_port, buffer_out_vector_0_44_port, 
      buffer_out_vector_0_43_port, buffer_out_vector_0_42_port, 
      buffer_out_vector_0_41_port, buffer_out_vector_0_40_port, 
      buffer_out_vector_0_39_port, buffer_out_vector_0_38_port, 
      buffer_out_vector_0_37_port, buffer_out_vector_0_36_port, 
      buffer_out_vector_0_35_port, buffer_out_vector_0_34_port, 
      buffer_out_vector_0_33_port, buffer_out_vector_0_32_port, 
      buffer_out_vector_0_31_port, buffer_out_vector_0_30_port, 
      buffer_out_vector_0_29_port, buffer_out_vector_0_28_port, 
      buffer_out_vector_0_27_port, buffer_out_vector_0_26_port, 
      buffer_out_vector_0_25_port, buffer_out_vector_0_24_port, 
      buffer_out_vector_0_23_port, buffer_out_vector_0_22_port, 
      buffer_out_vector_0_21_port, buffer_out_vector_0_20_port, 
      buffer_out_vector_0_19_port, buffer_out_vector_0_18_port, 
      buffer_out_vector_0_17_port, buffer_out_vector_0_16_port, 
      buffer_out_vector_0_15_port, buffer_out_vector_0_14_port, 
      buffer_out_vector_0_13_port, buffer_out_vector_0_12_port, 
      buffer_out_vector_0_11_port, buffer_out_vector_0_10_port, n1, n2, n3, n4,
      n5, n6, n7, n8 : std_logic;

begin
   header <= ( header_1_PACKET_LENGTH_3_port, header_1_PACKET_LENGTH_2_port, 
      header_1_PACKET_LENGTH_1_port, header_1_PACKET_LENGTH_0_port, 
      header_1_X_DEST_1_port, header_1_X_DEST_0_port, header_1_Y_DEST_1_port, 
      header_1_Y_DEST_0_port, header_1_Z_DEST_1_port, header_1_Z_DEST_0_port, 
      header_0_PACKET_LENGTH_3_port, header_0_PACKET_LENGTH_2_port, 
      header_0_PACKET_LENGTH_1_port, header_0_PACKET_LENGTH_0_port, 
      header_0_X_DEST_1_port, header_0_X_DEST_0_port, header_0_Y_DEST_1_port, 
      header_0_Y_DEST_0_port, header_0_Z_DEST_1_port, header_0_Z_DEST_0_port );
   
   U2 : AO22x1_ASAP7_75t_R port map( A1 => n3, A2 => 
                           buffer_out_vector_1_30_port, B1 => 
                           buffer_out_vector_0_30_port, B2 => n4, Y => 
                           data_transfer(30));
   U3 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_31_port, A2 => 
                           n3, B1 => buffer_out_vector_0_31_port, B2 => n4, Y 
                           => data_transfer(31));
   U4 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_32_port, A2 => 
                           n3, B1 => buffer_out_vector_0_32_port, B2 => n4, Y 
                           => data_transfer(32));
   U5 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_33_port, A2 => 
                           n3, B1 => buffer_out_vector_0_33_port, B2 => n4, Y 
                           => data_transfer(33));
   U6 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_34_port, A2 => 
                           n3, B1 => buffer_out_vector_0_34_port, B2 => n4, Y 
                           => data_transfer(34));
   U7 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_35_port, A2 => 
                           n3, B1 => buffer_out_vector_0_35_port, B2 => n6, Y 
                           => data_transfer(35));
   U8 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_36_port, A2 => 
                           n3, B1 => buffer_out_vector_0_36_port, B2 => n5, Y 
                           => data_transfer(36));
   U9 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_37_port, A2 => 
                           n3, B1 => buffer_out_vector_0_37_port, B2 => n7, Y 
                           => data_transfer(37));
   U10 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_38_port, A2 => 
                           n3, B1 => buffer_out_vector_0_38_port, B2 => n6, Y 
                           => data_transfer(38));
   U11 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_39_port, A2 => 
                           n3, B1 => buffer_out_vector_0_39_port, B2 => n5, Y 
                           => data_transfer(39));
   U12 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_40_port, A2 => 
                           n3, B1 => buffer_out_vector_0_40_port, B2 => n7, Y 
                           => data_transfer(40));
   U13 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_41_port, A2 => 
                           n3, B1 => buffer_out_vector_0_41_port, B2 => n6, Y 
                           => data_transfer(41));
   U14 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_42_port, A2 => 
                           n3, B1 => buffer_out_vector_0_42_port, B2 => n5, Y 
                           => data_transfer(42));
   U15 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_43_port, A2 => 
                           n3, B1 => buffer_out_vector_0_43_port, B2 => n7, Y 
                           => data_transfer(43));
   U16 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_44_port, A2 => 
                           n3, B1 => buffer_out_vector_0_44_port, B2 => n6, Y 
                           => data_transfer(44));
   U17 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_45_port, A2 => 
                           n3, B1 => buffer_out_vector_0_45_port, B2 => n5, Y 
                           => data_transfer(45));
   U18 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_46_port, A2 => 
                           n3, B1 => buffer_out_vector_0_46_port, B2 => n7, Y 
                           => data_transfer(46));
   U19 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_47_port, A2 => 
                           n3, B1 => buffer_out_vector_0_47_port, B2 => n7, Y 
                           => data_transfer(47));
   U20 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_48_port, A2 => 
                           n3, B1 => buffer_out_vector_0_48_port, B2 => n6, Y 
                           => data_transfer(48));
   U21 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_49_port, A2 => 
                           n3, B1 => buffer_out_vector_0_49_port, B2 => n5, Y 
                           => data_transfer(49));
   U22 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_50_port, A2 => 
                           n3, B1 => buffer_out_vector_0_50_port, B2 => n6, Y 
                           => data_transfer(50));
   U23 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_51_port, A2 => 
                           n2, B1 => buffer_out_vector_0_51_port, B2 => n7, Y 
                           => data_transfer(51));
   U24 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_52_port, A2 => 
                           n2, B1 => buffer_out_vector_0_52_port, B2 => n5, Y 
                           => data_transfer(52));
   U25 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_53_port, A2 => 
                           n2, B1 => buffer_out_vector_0_53_port, B2 => n6, Y 
                           => data_transfer(53));
   U26 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_54_port, A2 => 
                           n2, B1 => buffer_out_vector_0_54_port, B2 => n7, Y 
                           => data_transfer(54));
   U27 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_55_port, A2 => 
                           n2, B1 => buffer_out_vector_0_55_port, B2 => n5, Y 
                           => data_transfer(55));
   U28 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_56_port, A2 => 
                           n2, B1 => buffer_out_vector_0_56_port, B2 => n6, Y 
                           => data_transfer(56));
   U29 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_57_port, A2 => 
                           n2, B1 => buffer_out_vector_0_57_port, B2 => n7, Y 
                           => data_transfer(57));
   U30 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_58_port, A2 => 
                           n2, B1 => buffer_out_vector_0_58_port, B2 => n5, Y 
                           => data_transfer(58));
   U31 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_59_port, A2 => 
                           n2, B1 => buffer_out_vector_0_59_port, B2 => n7, Y 
                           => data_transfer(59));
   U32 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_60_port, A2 => 
                           n2, B1 => buffer_out_vector_0_60_port, B2 => n6, Y 
                           => data_transfer(60));
   U33 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_61_port, A2 => 
                           n2, B1 => buffer_out_vector_0_61_port, B2 => n7, Y 
                           => data_transfer(61));
   U34 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_62_port, A2 => 
                           n2, B1 => buffer_out_vector_0_62_port, B2 => n5, Y 
                           => data_transfer(62));
   U35 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_63_port, A2 => 
                           n2, B1 => buffer_out_vector_0_63_port, B2 => n6, Y 
                           => data_transfer(63));
   U36 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_0_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_0_port, B2 => n7
                           , Y => data_transfer(0));
   U37 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_1_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_1_port, B2 => n6
                           , Y => data_transfer(1));
   U38 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_2_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_2_port, B2 => n5
                           , Y => data_transfer(2));
   U39 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_3_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_3_port, B2 => n5
                           , Y => data_transfer(3));
   U40 : AO22x1_ASAP7_75t_R port map( A1 => header_1_X_DEST_0_port, A2 => n2, 
                           B1 => header_0_X_DEST_0_port, B2 => n5, Y => 
                           data_transfer(4));
   U41 : AO22x1_ASAP7_75t_R port map( A1 => header_1_X_DEST_1_port, A2 => n2, 
                           B1 => header_0_X_DEST_1_port, B2 => n5, Y => 
                           data_transfer(5));
   U42 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Y_DEST_0_port, A2 => n2, 
                           B1 => header_0_Y_DEST_0_port, B2 => n5, Y => 
                           data_transfer(6));
   U43 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Y_DEST_1_port, A2 => n2, 
                           B1 => header_0_Y_DEST_1_port, B2 => n5, Y => 
                           data_transfer(7));
   U44 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Z_DEST_0_port, A2 => n2, 
                           B1 => header_0_Z_DEST_0_port, B2 => n5, Y => 
                           data_transfer(8));
   U45 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Z_DEST_1_port, A2 => n2, 
                           B1 => header_0_Z_DEST_1_port, B2 => n5, Y => 
                           data_transfer(9));
   U46 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_10_port, A2 => 
                           n2, B1 => buffer_out_vector_0_10_port, B2 => n5, Y 
                           => data_transfer(10));
   U47 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_11_port, A2 => 
                           n2, B1 => buffer_out_vector_0_11_port, B2 => n6, Y 
                           => data_transfer(11));
   U48 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_12_port, A2 => 
                           n2, B1 => buffer_out_vector_0_12_port, B2 => n6, Y 
                           => data_transfer(12));
   U49 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_13_port, A2 => 
                           n2, B1 => buffer_out_vector_0_13_port, B2 => n6, Y 
                           => data_transfer(13));
   U50 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_14_port, A2 => 
                           n2, B1 => buffer_out_vector_0_14_port, B2 => n6, Y 
                           => data_transfer(14));
   U51 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_15_port, A2 => 
                           n2, B1 => buffer_out_vector_0_15_port, B2 => n6, Y 
                           => data_transfer(15));
   U52 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_16_port, A2 => 
                           n2, B1 => buffer_out_vector_0_16_port, B2 => n6, Y 
                           => data_transfer(16));
   U53 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_17_port, A2 => 
                           n2, B1 => buffer_out_vector_0_17_port, B2 => n6, Y 
                           => data_transfer(17));
   U54 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_18_port, A2 => 
                           n2, B1 => buffer_out_vector_0_18_port, B2 => n6, Y 
                           => data_transfer(18));
   U55 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_19_port, A2 => 
                           n2, B1 => buffer_out_vector_0_19_port, B2 => n7, Y 
                           => data_transfer(19));
   U56 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_20_port, A2 => 
                           n2, B1 => buffer_out_vector_0_20_port, B2 => n7, Y 
                           => data_transfer(20));
   U57 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_21_port, A2 => 
                           n2, B1 => buffer_out_vector_0_21_port, B2 => n7, Y 
                           => data_transfer(21));
   U58 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_22_port, A2 => 
                           n2, B1 => buffer_out_vector_0_22_port, B2 => n7, Y 
                           => data_transfer(22));
   U59 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_23_port, A2 => 
                           n2, B1 => buffer_out_vector_0_23_port, B2 => n7, Y 
                           => data_transfer(23));
   U60 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_24_port, A2 => 
                           n2, B1 => buffer_out_vector_0_24_port, B2 => n7, Y 
                           => data_transfer(24));
   U61 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_25_port, A2 => 
                           n2, B1 => buffer_out_vector_0_25_port, B2 => n7, Y 
                           => data_transfer(25));
   U62 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_26_port, A2 => 
                           n2, B1 => buffer_out_vector_0_26_port, B2 => n7, Y 
                           => data_transfer(26));
   U63 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_27_port, A2 => 
                           n2, B1 => buffer_out_vector_0_27_port, B2 => n6, Y 
                           => data_transfer(27));
   U64 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_28_port, A2 => 
                           n2, B1 => buffer_out_vector_0_28_port, B2 => n5, Y 
                           => data_transfer(28));
   U65 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_29_port, A2 => 
                           n2, B1 => buffer_out_vector_0_29_port, B2 => n5, Y 
                           => data_transfer(29));
   fifo_i_0 : fifo_buff_depth2_8 port map( data_in(63) => data_rx(63), 
                           data_in(62) => data_rx(62), data_in(61) => 
                           data_rx(61), data_in(60) => data_rx(60), data_in(59)
                           => data_rx(59), data_in(58) => data_rx(58), 
                           data_in(57) => data_rx(57), data_in(56) => 
                           data_rx(56), data_in(55) => data_rx(55), data_in(54)
                           => data_rx(54), data_in(53) => data_rx(53), 
                           data_in(52) => data_rx(52), data_in(51) => 
                           data_rx(51), data_in(50) => data_rx(50), data_in(49)
                           => data_rx(49), data_in(48) => data_rx(48), 
                           data_in(47) => data_rx(47), data_in(46) => 
                           data_rx(46), data_in(45) => data_rx(45), data_in(44)
                           => data_rx(44), data_in(43) => data_rx(43), 
                           data_in(42) => data_rx(42), data_in(41) => 
                           data_rx(41), data_in(40) => data_rx(40), data_in(39)
                           => data_rx(39), data_in(38) => data_rx(38), 
                           data_in(37) => data_rx(37), data_in(36) => 
                           data_rx(36), data_in(35) => data_rx(35), data_in(34)
                           => data_rx(34), data_in(33) => data_rx(33), 
                           data_in(32) => data_rx(32), data_in(31) => 
                           data_rx(31), data_in(30) => data_rx(30), data_in(29)
                           => data_rx(29), data_in(28) => data_rx(28), 
                           data_in(27) => data_rx(27), data_in(26) => 
                           data_rx(26), data_in(25) => data_rx(25), data_in(24)
                           => data_rx(24), data_in(23) => data_rx(23), 
                           data_in(22) => data_rx(22), data_in(21) => 
                           data_rx(21), data_in(20) => data_rx(20), data_in(19)
                           => data_rx(19), data_in(18) => data_rx(18), 
                           data_in(17) => data_rx(17), data_in(16) => 
                           data_rx(16), data_in(15) => data_rx(15), data_in(14)
                           => data_rx(14), data_in(13) => data_rx(13), 
                           data_in(12) => data_rx(12), data_in(11) => 
                           data_rx(11), data_in(10) => data_rx(10), data_in(9) 
                           => data_rx(9), data_in(8) => data_rx(8), data_in(7) 
                           => data_rx(7), data_in(6) => data_rx(6), data_in(5) 
                           => data_rx(5), data_in(4) => data_rx(4), data_in(3) 
                           => data_rx(3), data_in(2) => data_rx(2), data_in(1) 
                           => data_rx(1), data_in(0) => data_rx(0), write_en =>
                           vc_write_rx(0), read_en => vc_transfer(0), clk => 
                           clk, rst => n8, data_out(63) => 
                           buffer_out_vector_0_63_port, data_out(62) => 
                           buffer_out_vector_0_62_port, data_out(61) => 
                           buffer_out_vector_0_61_port, data_out(60) => 
                           buffer_out_vector_0_60_port, data_out(59) => 
                           buffer_out_vector_0_59_port, data_out(58) => 
                           buffer_out_vector_0_58_port, data_out(57) => 
                           buffer_out_vector_0_57_port, data_out(56) => 
                           buffer_out_vector_0_56_port, data_out(55) => 
                           buffer_out_vector_0_55_port, data_out(54) => 
                           buffer_out_vector_0_54_port, data_out(53) => 
                           buffer_out_vector_0_53_port, data_out(52) => 
                           buffer_out_vector_0_52_port, data_out(51) => 
                           buffer_out_vector_0_51_port, data_out(50) => 
                           buffer_out_vector_0_50_port, data_out(49) => 
                           buffer_out_vector_0_49_port, data_out(48) => 
                           buffer_out_vector_0_48_port, data_out(47) => 
                           buffer_out_vector_0_47_port, data_out(46) => 
                           buffer_out_vector_0_46_port, data_out(45) => 
                           buffer_out_vector_0_45_port, data_out(44) => 
                           buffer_out_vector_0_44_port, data_out(43) => 
                           buffer_out_vector_0_43_port, data_out(42) => 
                           buffer_out_vector_0_42_port, data_out(41) => 
                           buffer_out_vector_0_41_port, data_out(40) => 
                           buffer_out_vector_0_40_port, data_out(39) => 
                           buffer_out_vector_0_39_port, data_out(38) => 
                           buffer_out_vector_0_38_port, data_out(37) => 
                           buffer_out_vector_0_37_port, data_out(36) => 
                           buffer_out_vector_0_36_port, data_out(35) => 
                           buffer_out_vector_0_35_port, data_out(34) => 
                           buffer_out_vector_0_34_port, data_out(33) => 
                           buffer_out_vector_0_33_port, data_out(32) => 
                           buffer_out_vector_0_32_port, data_out(31) => 
                           buffer_out_vector_0_31_port, data_out(30) => 
                           buffer_out_vector_0_30_port, data_out(29) => 
                           buffer_out_vector_0_29_port, data_out(28) => 
                           buffer_out_vector_0_28_port, data_out(27) => 
                           buffer_out_vector_0_27_port, data_out(26) => 
                           buffer_out_vector_0_26_port, data_out(25) => 
                           buffer_out_vector_0_25_port, data_out(24) => 
                           buffer_out_vector_0_24_port, data_out(23) => 
                           buffer_out_vector_0_23_port, data_out(22) => 
                           buffer_out_vector_0_22_port, data_out(21) => 
                           buffer_out_vector_0_21_port, data_out(20) => 
                           buffer_out_vector_0_20_port, data_out(19) => 
                           buffer_out_vector_0_19_port, data_out(18) => 
                           buffer_out_vector_0_18_port, data_out(17) => 
                           buffer_out_vector_0_17_port, data_out(16) => 
                           buffer_out_vector_0_16_port, data_out(15) => 
                           buffer_out_vector_0_15_port, data_out(14) => 
                           buffer_out_vector_0_14_port, data_out(13) => 
                           buffer_out_vector_0_13_port, data_out(12) => 
                           buffer_out_vector_0_12_port, data_out(11) => 
                           buffer_out_vector_0_11_port, data_out(10) => 
                           buffer_out_vector_0_10_port, data_out(9) => 
                           header_0_Z_DEST_1_port, data_out(8) => 
                           header_0_Z_DEST_0_port, data_out(7) => 
                           header_0_Y_DEST_1_port, data_out(6) => 
                           header_0_Y_DEST_0_port, data_out(5) => 
                           header_0_X_DEST_1_port, data_out(4) => 
                           header_0_X_DEST_0_port, data_out(3) => 
                           header_0_PACKET_LENGTH_3_port, data_out(2) => 
                           header_0_PACKET_LENGTH_2_port, data_out(1) => 
                           header_0_PACKET_LENGTH_1_port, data_out(0) => 
                           header_0_PACKET_LENGTH_0_port, valid_data => 
                           valid_data_vc(0));
   fifo_i_1 : fifo_buff_depth2_7 port map( data_in(63) => data_rx(63), 
                           data_in(62) => data_rx(62), data_in(61) => 
                           data_rx(61), data_in(60) => data_rx(60), data_in(59)
                           => data_rx(59), data_in(58) => data_rx(58), 
                           data_in(57) => data_rx(57), data_in(56) => 
                           data_rx(56), data_in(55) => data_rx(55), data_in(54)
                           => data_rx(54), data_in(53) => data_rx(53), 
                           data_in(52) => data_rx(52), data_in(51) => 
                           data_rx(51), data_in(50) => data_rx(50), data_in(49)
                           => data_rx(49), data_in(48) => data_rx(48), 
                           data_in(47) => data_rx(47), data_in(46) => 
                           data_rx(46), data_in(45) => data_rx(45), data_in(44)
                           => data_rx(44), data_in(43) => data_rx(43), 
                           data_in(42) => data_rx(42), data_in(41) => 
                           data_rx(41), data_in(40) => data_rx(40), data_in(39)
                           => data_rx(39), data_in(38) => data_rx(38), 
                           data_in(37) => data_rx(37), data_in(36) => 
                           data_rx(36), data_in(35) => data_rx(35), data_in(34)
                           => data_rx(34), data_in(33) => data_rx(33), 
                           data_in(32) => data_rx(32), data_in(31) => 
                           data_rx(31), data_in(30) => data_rx(30), data_in(29)
                           => data_rx(29), data_in(28) => data_rx(28), 
                           data_in(27) => data_rx(27), data_in(26) => 
                           data_rx(26), data_in(25) => data_rx(25), data_in(24)
                           => data_rx(24), data_in(23) => data_rx(23), 
                           data_in(22) => data_rx(22), data_in(21) => 
                           data_rx(21), data_in(20) => data_rx(20), data_in(19)
                           => data_rx(19), data_in(18) => data_rx(18), 
                           data_in(17) => data_rx(17), data_in(16) => 
                           data_rx(16), data_in(15) => data_rx(15), data_in(14)
                           => data_rx(14), data_in(13) => data_rx(13), 
                           data_in(12) => data_rx(12), data_in(11) => 
                           data_rx(11), data_in(10) => data_rx(10), data_in(9) 
                           => data_rx(9), data_in(8) => data_rx(8), data_in(7) 
                           => data_rx(7), data_in(6) => data_rx(6), data_in(5) 
                           => data_rx(5), data_in(4) => data_rx(4), data_in(3) 
                           => data_rx(3), data_in(2) => data_rx(2), data_in(1) 
                           => data_rx(1), data_in(0) => data_rx(0), write_en =>
                           vc_write_rx(1), read_en => n2, clk => clk, rst => n8
                           , data_out(63) => buffer_out_vector_1_63_port, 
                           data_out(62) => buffer_out_vector_1_62_port, 
                           data_out(61) => buffer_out_vector_1_61_port, 
                           data_out(60) => buffer_out_vector_1_60_port, 
                           data_out(59) => buffer_out_vector_1_59_port, 
                           data_out(58) => buffer_out_vector_1_58_port, 
                           data_out(57) => buffer_out_vector_1_57_port, 
                           data_out(56) => buffer_out_vector_1_56_port, 
                           data_out(55) => buffer_out_vector_1_55_port, 
                           data_out(54) => buffer_out_vector_1_54_port, 
                           data_out(53) => buffer_out_vector_1_53_port, 
                           data_out(52) => buffer_out_vector_1_52_port, 
                           data_out(51) => buffer_out_vector_1_51_port, 
                           data_out(50) => buffer_out_vector_1_50_port, 
                           data_out(49) => buffer_out_vector_1_49_port, 
                           data_out(48) => buffer_out_vector_1_48_port, 
                           data_out(47) => buffer_out_vector_1_47_port, 
                           data_out(46) => buffer_out_vector_1_46_port, 
                           data_out(45) => buffer_out_vector_1_45_port, 
                           data_out(44) => buffer_out_vector_1_44_port, 
                           data_out(43) => buffer_out_vector_1_43_port, 
                           data_out(42) => buffer_out_vector_1_42_port, 
                           data_out(41) => buffer_out_vector_1_41_port, 
                           data_out(40) => buffer_out_vector_1_40_port, 
                           data_out(39) => buffer_out_vector_1_39_port, 
                           data_out(38) => buffer_out_vector_1_38_port, 
                           data_out(37) => buffer_out_vector_1_37_port, 
                           data_out(36) => buffer_out_vector_1_36_port, 
                           data_out(35) => buffer_out_vector_1_35_port, 
                           data_out(34) => buffer_out_vector_1_34_port, 
                           data_out(33) => buffer_out_vector_1_33_port, 
                           data_out(32) => buffer_out_vector_1_32_port, 
                           data_out(31) => buffer_out_vector_1_31_port, 
                           data_out(30) => buffer_out_vector_1_30_port, 
                           data_out(29) => buffer_out_vector_1_29_port, 
                           data_out(28) => buffer_out_vector_1_28_port, 
                           data_out(27) => buffer_out_vector_1_27_port, 
                           data_out(26) => buffer_out_vector_1_26_port, 
                           data_out(25) => buffer_out_vector_1_25_port, 
                           data_out(24) => buffer_out_vector_1_24_port, 
                           data_out(23) => buffer_out_vector_1_23_port, 
                           data_out(22) => buffer_out_vector_1_22_port, 
                           data_out(21) => buffer_out_vector_1_21_port, 
                           data_out(20) => buffer_out_vector_1_20_port, 
                           data_out(19) => buffer_out_vector_1_19_port, 
                           data_out(18) => buffer_out_vector_1_18_port, 
                           data_out(17) => buffer_out_vector_1_17_port, 
                           data_out(16) => buffer_out_vector_1_16_port, 
                           data_out(15) => buffer_out_vector_1_15_port, 
                           data_out(14) => buffer_out_vector_1_14_port, 
                           data_out(13) => buffer_out_vector_1_13_port, 
                           data_out(12) => buffer_out_vector_1_12_port, 
                           data_out(11) => buffer_out_vector_1_11_port, 
                           data_out(10) => buffer_out_vector_1_10_port, 
                           data_out(9) => header_1_Z_DEST_1_port, data_out(8) 
                           => header_1_Z_DEST_0_port, data_out(7) => 
                           header_1_Y_DEST_1_port, data_out(6) => 
                           header_1_Y_DEST_0_port, data_out(5) => 
                           header_1_X_DEST_1_port, data_out(4) => 
                           header_1_X_DEST_0_port, data_out(3) => 
                           header_1_PACKET_LENGTH_3_port, data_out(2) => 
                           header_1_PACKET_LENGTH_2_port, data_out(1) => 
                           header_1_PACKET_LENGTH_1_port, data_out(0) => 
                           header_1_PACKET_LENGTH_0_port, valid_data => 
                           valid_data_vc(1));
   U1 : INVx1_ASAP7_75t_R port map( A => n4, Y => n2);
   U66 : INVx1_ASAP7_75t_R port map( A => n4, Y => n3);
   U67 : INVx1_ASAP7_75t_R port map( A => n1, Y => n4);
   U68 : INVx1_ASAP7_75t_R port map( A => n1, Y => n5);
   U69 : INVx1_ASAP7_75t_R port map( A => n1, Y => n6);
   U70 : INVx1_ASAP7_75t_R port map( A => n1, Y => n7);
   U71 : HB1xp67_ASAP7_75t_R port map( A => vc_transfer(1), Y => n1);
   U72 : HB1xp67_ASAP7_75t_R port map( A => rst, Y => n8);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity vc_input_buffer_2_0000000200000002_3 is

   port( clk, rst : in std_logic;  data_rx : in std_logic_vector (63 downto 0);
         vc_write_rx, vc_transfer : in std_logic_vector (1 downto 0);  
         valid_data_vc : out std_logic_vector (1 downto 0);  data_transfer : 
         out std_logic_vector (63 downto 0);  header : out std_logic_vector (19
         downto 0));

end vc_input_buffer_2_0000000200000002_3;

architecture SYN_rtl of vc_input_buffer_2_0000000200000002_3 is

   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component fifo_buff_depth2_5
      port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, 
            clk, rst : in std_logic;  data_out : out std_logic_vector (63 
            downto 0);  valid_data : out std_logic);
   end component;
   
   component fifo_buff_depth2_6
      port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, 
            clk, rst : in std_logic;  data_out : out std_logic_vector (63 
            downto 0);  valid_data : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal header_1_PACKET_LENGTH_3_port, header_1_PACKET_LENGTH_2_port, 
      header_1_PACKET_LENGTH_1_port, header_1_PACKET_LENGTH_0_port, 
      header_1_X_DEST_1_port, header_1_X_DEST_0_port, header_1_Y_DEST_1_port, 
      header_1_Y_DEST_0_port, header_1_Z_DEST_1_port, header_1_Z_DEST_0_port, 
      header_0_PACKET_LENGTH_3_port, header_0_PACKET_LENGTH_2_port, 
      header_0_PACKET_LENGTH_1_port, header_0_PACKET_LENGTH_0_port, 
      header_0_X_DEST_1_port, header_0_X_DEST_0_port, header_0_Y_DEST_1_port, 
      header_0_Y_DEST_0_port, header_0_Z_DEST_1_port, header_0_Z_DEST_0_port, 
      buffer_out_vector_1_63_port, buffer_out_vector_1_62_port, 
      buffer_out_vector_1_61_port, buffer_out_vector_1_60_port, 
      buffer_out_vector_1_59_port, buffer_out_vector_1_58_port, 
      buffer_out_vector_1_57_port, buffer_out_vector_1_56_port, 
      buffer_out_vector_1_55_port, buffer_out_vector_1_54_port, 
      buffer_out_vector_1_53_port, buffer_out_vector_1_52_port, 
      buffer_out_vector_1_51_port, buffer_out_vector_1_50_port, 
      buffer_out_vector_1_49_port, buffer_out_vector_1_48_port, 
      buffer_out_vector_1_47_port, buffer_out_vector_1_46_port, 
      buffer_out_vector_1_45_port, buffer_out_vector_1_44_port, 
      buffer_out_vector_1_43_port, buffer_out_vector_1_42_port, 
      buffer_out_vector_1_41_port, buffer_out_vector_1_40_port, 
      buffer_out_vector_1_39_port, buffer_out_vector_1_38_port, 
      buffer_out_vector_1_37_port, buffer_out_vector_1_36_port, 
      buffer_out_vector_1_35_port, buffer_out_vector_1_34_port, 
      buffer_out_vector_1_33_port, buffer_out_vector_1_32_port, 
      buffer_out_vector_1_31_port, buffer_out_vector_1_30_port, 
      buffer_out_vector_1_29_port, buffer_out_vector_1_28_port, 
      buffer_out_vector_1_27_port, buffer_out_vector_1_26_port, 
      buffer_out_vector_1_25_port, buffer_out_vector_1_24_port, 
      buffer_out_vector_1_23_port, buffer_out_vector_1_22_port, 
      buffer_out_vector_1_21_port, buffer_out_vector_1_20_port, 
      buffer_out_vector_1_19_port, buffer_out_vector_1_18_port, 
      buffer_out_vector_1_17_port, buffer_out_vector_1_16_port, 
      buffer_out_vector_1_15_port, buffer_out_vector_1_14_port, 
      buffer_out_vector_1_13_port, buffer_out_vector_1_12_port, 
      buffer_out_vector_1_11_port, buffer_out_vector_1_10_port, 
      buffer_out_vector_0_63_port, buffer_out_vector_0_62_port, 
      buffer_out_vector_0_61_port, buffer_out_vector_0_60_port, 
      buffer_out_vector_0_59_port, buffer_out_vector_0_58_port, 
      buffer_out_vector_0_57_port, buffer_out_vector_0_56_port, 
      buffer_out_vector_0_55_port, buffer_out_vector_0_54_port, 
      buffer_out_vector_0_53_port, buffer_out_vector_0_52_port, 
      buffer_out_vector_0_51_port, buffer_out_vector_0_50_port, 
      buffer_out_vector_0_49_port, buffer_out_vector_0_48_port, 
      buffer_out_vector_0_47_port, buffer_out_vector_0_46_port, 
      buffer_out_vector_0_45_port, buffer_out_vector_0_44_port, 
      buffer_out_vector_0_43_port, buffer_out_vector_0_42_port, 
      buffer_out_vector_0_41_port, buffer_out_vector_0_40_port, 
      buffer_out_vector_0_39_port, buffer_out_vector_0_38_port, 
      buffer_out_vector_0_37_port, buffer_out_vector_0_36_port, 
      buffer_out_vector_0_35_port, buffer_out_vector_0_34_port, 
      buffer_out_vector_0_33_port, buffer_out_vector_0_32_port, 
      buffer_out_vector_0_31_port, buffer_out_vector_0_30_port, 
      buffer_out_vector_0_29_port, buffer_out_vector_0_28_port, 
      buffer_out_vector_0_27_port, buffer_out_vector_0_26_port, 
      buffer_out_vector_0_25_port, buffer_out_vector_0_24_port, 
      buffer_out_vector_0_23_port, buffer_out_vector_0_22_port, 
      buffer_out_vector_0_21_port, buffer_out_vector_0_20_port, 
      buffer_out_vector_0_19_port, buffer_out_vector_0_18_port, 
      buffer_out_vector_0_17_port, buffer_out_vector_0_16_port, 
      buffer_out_vector_0_15_port, buffer_out_vector_0_14_port, 
      buffer_out_vector_0_13_port, buffer_out_vector_0_12_port, 
      buffer_out_vector_0_11_port, buffer_out_vector_0_10_port, n1, n2, n3, n4,
      n5, n6, n7, n8 : std_logic;

begin
   header <= ( header_1_PACKET_LENGTH_3_port, header_1_PACKET_LENGTH_2_port, 
      header_1_PACKET_LENGTH_1_port, header_1_PACKET_LENGTH_0_port, 
      header_1_X_DEST_1_port, header_1_X_DEST_0_port, header_1_Y_DEST_1_port, 
      header_1_Y_DEST_0_port, header_1_Z_DEST_1_port, header_1_Z_DEST_0_port, 
      header_0_PACKET_LENGTH_3_port, header_0_PACKET_LENGTH_2_port, 
      header_0_PACKET_LENGTH_1_port, header_0_PACKET_LENGTH_0_port, 
      header_0_X_DEST_1_port, header_0_X_DEST_0_port, header_0_Y_DEST_1_port, 
      header_0_Y_DEST_0_port, header_0_Z_DEST_1_port, header_0_Z_DEST_0_port );
   
   U2 : AO22x1_ASAP7_75t_R port map( A1 => n3, A2 => 
                           buffer_out_vector_1_30_port, B1 => 
                           buffer_out_vector_0_30_port, B2 => n4, Y => 
                           data_transfer(30));
   U3 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_31_port, A2 => 
                           n3, B1 => buffer_out_vector_0_31_port, B2 => n4, Y 
                           => data_transfer(31));
   U4 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_32_port, A2 => 
                           n3, B1 => buffer_out_vector_0_32_port, B2 => n4, Y 
                           => data_transfer(32));
   U5 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_33_port, A2 => 
                           n3, B1 => buffer_out_vector_0_33_port, B2 => n4, Y 
                           => data_transfer(33));
   U6 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_34_port, A2 => 
                           n3, B1 => buffer_out_vector_0_34_port, B2 => n4, Y 
                           => data_transfer(34));
   U7 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_35_port, A2 => 
                           n3, B1 => buffer_out_vector_0_35_port, B2 => n6, Y 
                           => data_transfer(35));
   U8 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_36_port, A2 => 
                           n3, B1 => buffer_out_vector_0_36_port, B2 => n5, Y 
                           => data_transfer(36));
   U9 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_37_port, A2 => 
                           n3, B1 => buffer_out_vector_0_37_port, B2 => n7, Y 
                           => data_transfer(37));
   U10 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_38_port, A2 => 
                           n3, B1 => buffer_out_vector_0_38_port, B2 => n6, Y 
                           => data_transfer(38));
   U11 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_39_port, A2 => 
                           n3, B1 => buffer_out_vector_0_39_port, B2 => n5, Y 
                           => data_transfer(39));
   U12 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_40_port, A2 => 
                           n3, B1 => buffer_out_vector_0_40_port, B2 => n7, Y 
                           => data_transfer(40));
   U13 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_41_port, A2 => 
                           n3, B1 => buffer_out_vector_0_41_port, B2 => n6, Y 
                           => data_transfer(41));
   U14 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_42_port, A2 => 
                           n3, B1 => buffer_out_vector_0_42_port, B2 => n5, Y 
                           => data_transfer(42));
   U15 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_43_port, A2 => 
                           n3, B1 => buffer_out_vector_0_43_port, B2 => n7, Y 
                           => data_transfer(43));
   U16 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_44_port, A2 => 
                           n3, B1 => buffer_out_vector_0_44_port, B2 => n7, Y 
                           => data_transfer(44));
   U17 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_45_port, A2 => 
                           n3, B1 => buffer_out_vector_0_45_port, B2 => n6, Y 
                           => data_transfer(45));
   U18 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_46_port, A2 => 
                           n3, B1 => buffer_out_vector_0_46_port, B2 => n5, Y 
                           => data_transfer(46));
   U19 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_47_port, A2 => 
                           n3, B1 => buffer_out_vector_0_47_port, B2 => n6, Y 
                           => data_transfer(47));
   U20 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_48_port, A2 => 
                           n3, B1 => buffer_out_vector_0_48_port, B2 => n6, Y 
                           => data_transfer(48));
   U21 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_49_port, A2 => 
                           n3, B1 => buffer_out_vector_0_49_port, B2 => n7, Y 
                           => data_transfer(49));
   U22 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_50_port, A2 => 
                           n3, B1 => buffer_out_vector_0_50_port, B2 => n6, Y 
                           => data_transfer(50));
   U23 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_51_port, A2 => 
                           n2, B1 => buffer_out_vector_0_51_port, B2 => n7, Y 
                           => data_transfer(51));
   U24 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_52_port, A2 => 
                           n2, B1 => buffer_out_vector_0_52_port, B2 => n5, Y 
                           => data_transfer(52));
   U25 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_53_port, A2 => 
                           n2, B1 => buffer_out_vector_0_53_port, B2 => n5, Y 
                           => data_transfer(53));
   U26 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_54_port, A2 => 
                           n2, B1 => buffer_out_vector_0_54_port, B2 => n7, Y 
                           => data_transfer(54));
   U27 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_55_port, A2 => 
                           n2, B1 => buffer_out_vector_0_55_port, B2 => n6, Y 
                           => data_transfer(55));
   U28 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_56_port, A2 => 
                           n2, B1 => buffer_out_vector_0_56_port, B2 => n7, Y 
                           => data_transfer(56));
   U29 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_57_port, A2 => 
                           n2, B1 => buffer_out_vector_0_57_port, B2 => n7, Y 
                           => data_transfer(57));
   U30 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_58_port, A2 => 
                           n2, B1 => buffer_out_vector_0_58_port, B2 => n6, Y 
                           => data_transfer(58));
   U31 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_59_port, A2 => 
                           n2, B1 => buffer_out_vector_0_59_port, B2 => n5, Y 
                           => data_transfer(59));
   U32 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_60_port, A2 => 
                           n2, B1 => buffer_out_vector_0_60_port, B2 => n6, Y 
                           => data_transfer(60));
   U33 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_61_port, A2 => 
                           n2, B1 => buffer_out_vector_0_61_port, B2 => n6, Y 
                           => data_transfer(61));
   U34 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_62_port, A2 => 
                           n2, B1 => buffer_out_vector_0_62_port, B2 => n7, Y 
                           => data_transfer(62));
   U35 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_63_port, A2 => 
                           n2, B1 => buffer_out_vector_0_63_port, B2 => n5, Y 
                           => data_transfer(63));
   U36 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_0_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_0_port, B2 => n7
                           , Y => data_transfer(0));
   U37 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_1_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_1_port, B2 => n6
                           , Y => data_transfer(1));
   U38 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_2_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_2_port, B2 => n5
                           , Y => data_transfer(2));
   U39 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_3_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_3_port, B2 => n5
                           , Y => data_transfer(3));
   U40 : AO22x1_ASAP7_75t_R port map( A1 => header_1_X_DEST_0_port, A2 => n2, 
                           B1 => header_0_X_DEST_0_port, B2 => n5, Y => 
                           data_transfer(4));
   U41 : AO22x1_ASAP7_75t_R port map( A1 => header_1_X_DEST_1_port, A2 => n2, 
                           B1 => header_0_X_DEST_1_port, B2 => n5, Y => 
                           data_transfer(5));
   U42 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Y_DEST_0_port, A2 => n2, 
                           B1 => header_0_Y_DEST_0_port, B2 => n5, Y => 
                           data_transfer(6));
   U43 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Y_DEST_1_port, A2 => n2, 
                           B1 => header_0_Y_DEST_1_port, B2 => n5, Y => 
                           data_transfer(7));
   U44 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Z_DEST_0_port, A2 => n2, 
                           B1 => header_0_Z_DEST_0_port, B2 => n5, Y => 
                           data_transfer(8));
   U45 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Z_DEST_1_port, A2 => n2, 
                           B1 => header_0_Z_DEST_1_port, B2 => n5, Y => 
                           data_transfer(9));
   U46 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_10_port, A2 => 
                           n2, B1 => buffer_out_vector_0_10_port, B2 => n5, Y 
                           => data_transfer(10));
   U47 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_11_port, A2 => 
                           n2, B1 => buffer_out_vector_0_11_port, B2 => n6, Y 
                           => data_transfer(11));
   U48 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_12_port, A2 => 
                           n2, B1 => buffer_out_vector_0_12_port, B2 => n6, Y 
                           => data_transfer(12));
   U49 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_13_port, A2 => 
                           n2, B1 => buffer_out_vector_0_13_port, B2 => n6, Y 
                           => data_transfer(13));
   U50 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_14_port, A2 => 
                           n2, B1 => buffer_out_vector_0_14_port, B2 => n6, Y 
                           => data_transfer(14));
   U51 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_15_port, A2 => 
                           n2, B1 => buffer_out_vector_0_15_port, B2 => n6, Y 
                           => data_transfer(15));
   U52 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_16_port, A2 => 
                           n2, B1 => buffer_out_vector_0_16_port, B2 => n6, Y 
                           => data_transfer(16));
   U53 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_17_port, A2 => 
                           n2, B1 => buffer_out_vector_0_17_port, B2 => n6, Y 
                           => data_transfer(17));
   U54 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_18_port, A2 => 
                           n2, B1 => buffer_out_vector_0_18_port, B2 => n6, Y 
                           => data_transfer(18));
   U55 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_19_port, A2 => 
                           n2, B1 => buffer_out_vector_0_19_port, B2 => n7, Y 
                           => data_transfer(19));
   U56 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_20_port, A2 => 
                           n2, B1 => buffer_out_vector_0_20_port, B2 => n7, Y 
                           => data_transfer(20));
   U57 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_21_port, A2 => 
                           n2, B1 => buffer_out_vector_0_21_port, B2 => n7, Y 
                           => data_transfer(21));
   U58 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_22_port, A2 => 
                           n2, B1 => buffer_out_vector_0_22_port, B2 => n7, Y 
                           => data_transfer(22));
   U59 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_23_port, A2 => 
                           n2, B1 => buffer_out_vector_0_23_port, B2 => n7, Y 
                           => data_transfer(23));
   U60 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_24_port, A2 => 
                           n2, B1 => buffer_out_vector_0_24_port, B2 => n7, Y 
                           => data_transfer(24));
   U61 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_25_port, A2 => 
                           n2, B1 => buffer_out_vector_0_25_port, B2 => n7, Y 
                           => data_transfer(25));
   U62 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_26_port, A2 => 
                           n2, B1 => buffer_out_vector_0_26_port, B2 => n7, Y 
                           => data_transfer(26));
   U63 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_27_port, A2 => 
                           n2, B1 => buffer_out_vector_0_27_port, B2 => n5, Y 
                           => data_transfer(27));
   U64 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_28_port, A2 => 
                           n2, B1 => buffer_out_vector_0_28_port, B2 => n5, Y 
                           => data_transfer(28));
   U65 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_29_port, A2 => 
                           n2, B1 => buffer_out_vector_0_29_port, B2 => n5, Y 
                           => data_transfer(29));
   fifo_i_0 : fifo_buff_depth2_6 port map( data_in(63) => data_rx(63), 
                           data_in(62) => data_rx(62), data_in(61) => 
                           data_rx(61), data_in(60) => data_rx(60), data_in(59)
                           => data_rx(59), data_in(58) => data_rx(58), 
                           data_in(57) => data_rx(57), data_in(56) => 
                           data_rx(56), data_in(55) => data_rx(55), data_in(54)
                           => data_rx(54), data_in(53) => data_rx(53), 
                           data_in(52) => data_rx(52), data_in(51) => 
                           data_rx(51), data_in(50) => data_rx(50), data_in(49)
                           => data_rx(49), data_in(48) => data_rx(48), 
                           data_in(47) => data_rx(47), data_in(46) => 
                           data_rx(46), data_in(45) => data_rx(45), data_in(44)
                           => data_rx(44), data_in(43) => data_rx(43), 
                           data_in(42) => data_rx(42), data_in(41) => 
                           data_rx(41), data_in(40) => data_rx(40), data_in(39)
                           => data_rx(39), data_in(38) => data_rx(38), 
                           data_in(37) => data_rx(37), data_in(36) => 
                           data_rx(36), data_in(35) => data_rx(35), data_in(34)
                           => data_rx(34), data_in(33) => data_rx(33), 
                           data_in(32) => data_rx(32), data_in(31) => 
                           data_rx(31), data_in(30) => data_rx(30), data_in(29)
                           => data_rx(29), data_in(28) => data_rx(28), 
                           data_in(27) => data_rx(27), data_in(26) => 
                           data_rx(26), data_in(25) => data_rx(25), data_in(24)
                           => data_rx(24), data_in(23) => data_rx(23), 
                           data_in(22) => data_rx(22), data_in(21) => 
                           data_rx(21), data_in(20) => data_rx(20), data_in(19)
                           => data_rx(19), data_in(18) => data_rx(18), 
                           data_in(17) => data_rx(17), data_in(16) => 
                           data_rx(16), data_in(15) => data_rx(15), data_in(14)
                           => data_rx(14), data_in(13) => data_rx(13), 
                           data_in(12) => data_rx(12), data_in(11) => 
                           data_rx(11), data_in(10) => data_rx(10), data_in(9) 
                           => data_rx(9), data_in(8) => data_rx(8), data_in(7) 
                           => data_rx(7), data_in(6) => data_rx(6), data_in(5) 
                           => data_rx(5), data_in(4) => data_rx(4), data_in(3) 
                           => data_rx(3), data_in(2) => data_rx(2), data_in(1) 
                           => data_rx(1), data_in(0) => data_rx(0), write_en =>
                           vc_write_rx(0), read_en => vc_transfer(0), clk => 
                           clk, rst => n8, data_out(63) => 
                           buffer_out_vector_0_63_port, data_out(62) => 
                           buffer_out_vector_0_62_port, data_out(61) => 
                           buffer_out_vector_0_61_port, data_out(60) => 
                           buffer_out_vector_0_60_port, data_out(59) => 
                           buffer_out_vector_0_59_port, data_out(58) => 
                           buffer_out_vector_0_58_port, data_out(57) => 
                           buffer_out_vector_0_57_port, data_out(56) => 
                           buffer_out_vector_0_56_port, data_out(55) => 
                           buffer_out_vector_0_55_port, data_out(54) => 
                           buffer_out_vector_0_54_port, data_out(53) => 
                           buffer_out_vector_0_53_port, data_out(52) => 
                           buffer_out_vector_0_52_port, data_out(51) => 
                           buffer_out_vector_0_51_port, data_out(50) => 
                           buffer_out_vector_0_50_port, data_out(49) => 
                           buffer_out_vector_0_49_port, data_out(48) => 
                           buffer_out_vector_0_48_port, data_out(47) => 
                           buffer_out_vector_0_47_port, data_out(46) => 
                           buffer_out_vector_0_46_port, data_out(45) => 
                           buffer_out_vector_0_45_port, data_out(44) => 
                           buffer_out_vector_0_44_port, data_out(43) => 
                           buffer_out_vector_0_43_port, data_out(42) => 
                           buffer_out_vector_0_42_port, data_out(41) => 
                           buffer_out_vector_0_41_port, data_out(40) => 
                           buffer_out_vector_0_40_port, data_out(39) => 
                           buffer_out_vector_0_39_port, data_out(38) => 
                           buffer_out_vector_0_38_port, data_out(37) => 
                           buffer_out_vector_0_37_port, data_out(36) => 
                           buffer_out_vector_0_36_port, data_out(35) => 
                           buffer_out_vector_0_35_port, data_out(34) => 
                           buffer_out_vector_0_34_port, data_out(33) => 
                           buffer_out_vector_0_33_port, data_out(32) => 
                           buffer_out_vector_0_32_port, data_out(31) => 
                           buffer_out_vector_0_31_port, data_out(30) => 
                           buffer_out_vector_0_30_port, data_out(29) => 
                           buffer_out_vector_0_29_port, data_out(28) => 
                           buffer_out_vector_0_28_port, data_out(27) => 
                           buffer_out_vector_0_27_port, data_out(26) => 
                           buffer_out_vector_0_26_port, data_out(25) => 
                           buffer_out_vector_0_25_port, data_out(24) => 
                           buffer_out_vector_0_24_port, data_out(23) => 
                           buffer_out_vector_0_23_port, data_out(22) => 
                           buffer_out_vector_0_22_port, data_out(21) => 
                           buffer_out_vector_0_21_port, data_out(20) => 
                           buffer_out_vector_0_20_port, data_out(19) => 
                           buffer_out_vector_0_19_port, data_out(18) => 
                           buffer_out_vector_0_18_port, data_out(17) => 
                           buffer_out_vector_0_17_port, data_out(16) => 
                           buffer_out_vector_0_16_port, data_out(15) => 
                           buffer_out_vector_0_15_port, data_out(14) => 
                           buffer_out_vector_0_14_port, data_out(13) => 
                           buffer_out_vector_0_13_port, data_out(12) => 
                           buffer_out_vector_0_12_port, data_out(11) => 
                           buffer_out_vector_0_11_port, data_out(10) => 
                           buffer_out_vector_0_10_port, data_out(9) => 
                           header_0_Z_DEST_1_port, data_out(8) => 
                           header_0_Z_DEST_0_port, data_out(7) => 
                           header_0_Y_DEST_1_port, data_out(6) => 
                           header_0_Y_DEST_0_port, data_out(5) => 
                           header_0_X_DEST_1_port, data_out(4) => 
                           header_0_X_DEST_0_port, data_out(3) => 
                           header_0_PACKET_LENGTH_3_port, data_out(2) => 
                           header_0_PACKET_LENGTH_2_port, data_out(1) => 
                           header_0_PACKET_LENGTH_1_port, data_out(0) => 
                           header_0_PACKET_LENGTH_0_port, valid_data => 
                           valid_data_vc(0));
   fifo_i_1 : fifo_buff_depth2_5 port map( data_in(63) => data_rx(63), 
                           data_in(62) => data_rx(62), data_in(61) => 
                           data_rx(61), data_in(60) => data_rx(60), data_in(59)
                           => data_rx(59), data_in(58) => data_rx(58), 
                           data_in(57) => data_rx(57), data_in(56) => 
                           data_rx(56), data_in(55) => data_rx(55), data_in(54)
                           => data_rx(54), data_in(53) => data_rx(53), 
                           data_in(52) => data_rx(52), data_in(51) => 
                           data_rx(51), data_in(50) => data_rx(50), data_in(49)
                           => data_rx(49), data_in(48) => data_rx(48), 
                           data_in(47) => data_rx(47), data_in(46) => 
                           data_rx(46), data_in(45) => data_rx(45), data_in(44)
                           => data_rx(44), data_in(43) => data_rx(43), 
                           data_in(42) => data_rx(42), data_in(41) => 
                           data_rx(41), data_in(40) => data_rx(40), data_in(39)
                           => data_rx(39), data_in(38) => data_rx(38), 
                           data_in(37) => data_rx(37), data_in(36) => 
                           data_rx(36), data_in(35) => data_rx(35), data_in(34)
                           => data_rx(34), data_in(33) => data_rx(33), 
                           data_in(32) => data_rx(32), data_in(31) => 
                           data_rx(31), data_in(30) => data_rx(30), data_in(29)
                           => data_rx(29), data_in(28) => data_rx(28), 
                           data_in(27) => data_rx(27), data_in(26) => 
                           data_rx(26), data_in(25) => data_rx(25), data_in(24)
                           => data_rx(24), data_in(23) => data_rx(23), 
                           data_in(22) => data_rx(22), data_in(21) => 
                           data_rx(21), data_in(20) => data_rx(20), data_in(19)
                           => data_rx(19), data_in(18) => data_rx(18), 
                           data_in(17) => data_rx(17), data_in(16) => 
                           data_rx(16), data_in(15) => data_rx(15), data_in(14)
                           => data_rx(14), data_in(13) => data_rx(13), 
                           data_in(12) => data_rx(12), data_in(11) => 
                           data_rx(11), data_in(10) => data_rx(10), data_in(9) 
                           => data_rx(9), data_in(8) => data_rx(8), data_in(7) 
                           => data_rx(7), data_in(6) => data_rx(6), data_in(5) 
                           => data_rx(5), data_in(4) => data_rx(4), data_in(3) 
                           => data_rx(3), data_in(2) => data_rx(2), data_in(1) 
                           => data_rx(1), data_in(0) => data_rx(0), write_en =>
                           vc_write_rx(1), read_en => n2, clk => clk, rst => n8
                           , data_out(63) => buffer_out_vector_1_63_port, 
                           data_out(62) => buffer_out_vector_1_62_port, 
                           data_out(61) => buffer_out_vector_1_61_port, 
                           data_out(60) => buffer_out_vector_1_60_port, 
                           data_out(59) => buffer_out_vector_1_59_port, 
                           data_out(58) => buffer_out_vector_1_58_port, 
                           data_out(57) => buffer_out_vector_1_57_port, 
                           data_out(56) => buffer_out_vector_1_56_port, 
                           data_out(55) => buffer_out_vector_1_55_port, 
                           data_out(54) => buffer_out_vector_1_54_port, 
                           data_out(53) => buffer_out_vector_1_53_port, 
                           data_out(52) => buffer_out_vector_1_52_port, 
                           data_out(51) => buffer_out_vector_1_51_port, 
                           data_out(50) => buffer_out_vector_1_50_port, 
                           data_out(49) => buffer_out_vector_1_49_port, 
                           data_out(48) => buffer_out_vector_1_48_port, 
                           data_out(47) => buffer_out_vector_1_47_port, 
                           data_out(46) => buffer_out_vector_1_46_port, 
                           data_out(45) => buffer_out_vector_1_45_port, 
                           data_out(44) => buffer_out_vector_1_44_port, 
                           data_out(43) => buffer_out_vector_1_43_port, 
                           data_out(42) => buffer_out_vector_1_42_port, 
                           data_out(41) => buffer_out_vector_1_41_port, 
                           data_out(40) => buffer_out_vector_1_40_port, 
                           data_out(39) => buffer_out_vector_1_39_port, 
                           data_out(38) => buffer_out_vector_1_38_port, 
                           data_out(37) => buffer_out_vector_1_37_port, 
                           data_out(36) => buffer_out_vector_1_36_port, 
                           data_out(35) => buffer_out_vector_1_35_port, 
                           data_out(34) => buffer_out_vector_1_34_port, 
                           data_out(33) => buffer_out_vector_1_33_port, 
                           data_out(32) => buffer_out_vector_1_32_port, 
                           data_out(31) => buffer_out_vector_1_31_port, 
                           data_out(30) => buffer_out_vector_1_30_port, 
                           data_out(29) => buffer_out_vector_1_29_port, 
                           data_out(28) => buffer_out_vector_1_28_port, 
                           data_out(27) => buffer_out_vector_1_27_port, 
                           data_out(26) => buffer_out_vector_1_26_port, 
                           data_out(25) => buffer_out_vector_1_25_port, 
                           data_out(24) => buffer_out_vector_1_24_port, 
                           data_out(23) => buffer_out_vector_1_23_port, 
                           data_out(22) => buffer_out_vector_1_22_port, 
                           data_out(21) => buffer_out_vector_1_21_port, 
                           data_out(20) => buffer_out_vector_1_20_port, 
                           data_out(19) => buffer_out_vector_1_19_port, 
                           data_out(18) => buffer_out_vector_1_18_port, 
                           data_out(17) => buffer_out_vector_1_17_port, 
                           data_out(16) => buffer_out_vector_1_16_port, 
                           data_out(15) => buffer_out_vector_1_15_port, 
                           data_out(14) => buffer_out_vector_1_14_port, 
                           data_out(13) => buffer_out_vector_1_13_port, 
                           data_out(12) => buffer_out_vector_1_12_port, 
                           data_out(11) => buffer_out_vector_1_11_port, 
                           data_out(10) => buffer_out_vector_1_10_port, 
                           data_out(9) => header_1_Z_DEST_1_port, data_out(8) 
                           => header_1_Z_DEST_0_port, data_out(7) => 
                           header_1_Y_DEST_1_port, data_out(6) => 
                           header_1_Y_DEST_0_port, data_out(5) => 
                           header_1_X_DEST_1_port, data_out(4) => 
                           header_1_X_DEST_0_port, data_out(3) => 
                           header_1_PACKET_LENGTH_3_port, data_out(2) => 
                           header_1_PACKET_LENGTH_2_port, data_out(1) => 
                           header_1_PACKET_LENGTH_1_port, data_out(0) => 
                           header_1_PACKET_LENGTH_0_port, valid_data => 
                           valid_data_vc(1));
   U1 : INVx1_ASAP7_75t_R port map( A => n4, Y => n2);
   U66 : INVx1_ASAP7_75t_R port map( A => n4, Y => n3);
   U67 : INVx1_ASAP7_75t_R port map( A => n1, Y => n4);
   U68 : INVx1_ASAP7_75t_R port map( A => n1, Y => n5);
   U69 : INVx1_ASAP7_75t_R port map( A => n1, Y => n6);
   U70 : INVx1_ASAP7_75t_R port map( A => n1, Y => n7);
   U71 : HB1xp67_ASAP7_75t_R port map( A => vc_transfer(1), Y => n1);
   U72 : HB1xp67_ASAP7_75t_R port map( A => rst, Y => n8);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity vc_input_buffer_2_0000000200000002_2 is

   port( clk, rst : in std_logic;  data_rx : in std_logic_vector (63 downto 0);
         vc_write_rx, vc_transfer : in std_logic_vector (1 downto 0);  
         valid_data_vc : out std_logic_vector (1 downto 0);  data_transfer : 
         out std_logic_vector (63 downto 0);  header : out std_logic_vector (19
         downto 0));

end vc_input_buffer_2_0000000200000002_2;

architecture SYN_rtl of vc_input_buffer_2_0000000200000002_2 is

   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component fifo_buff_depth2_3
      port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, 
            clk, rst : in std_logic;  data_out : out std_logic_vector (63 
            downto 0);  valid_data : out std_logic);
   end component;
   
   component fifo_buff_depth2_4
      port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, 
            clk, rst : in std_logic;  data_out : out std_logic_vector (63 
            downto 0);  valid_data : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal header_1_PACKET_LENGTH_3_port, header_1_PACKET_LENGTH_2_port, 
      header_1_PACKET_LENGTH_1_port, header_1_PACKET_LENGTH_0_port, 
      header_1_X_DEST_1_port, header_1_X_DEST_0_port, header_1_Y_DEST_1_port, 
      header_1_Y_DEST_0_port, header_1_Z_DEST_1_port, header_1_Z_DEST_0_port, 
      header_0_PACKET_LENGTH_3_port, header_0_PACKET_LENGTH_2_port, 
      header_0_PACKET_LENGTH_1_port, header_0_PACKET_LENGTH_0_port, 
      header_0_X_DEST_1_port, header_0_X_DEST_0_port, header_0_Y_DEST_1_port, 
      header_0_Y_DEST_0_port, header_0_Z_DEST_1_port, header_0_Z_DEST_0_port, 
      buffer_out_vector_1_63_port, buffer_out_vector_1_62_port, 
      buffer_out_vector_1_61_port, buffer_out_vector_1_60_port, 
      buffer_out_vector_1_59_port, buffer_out_vector_1_58_port, 
      buffer_out_vector_1_57_port, buffer_out_vector_1_56_port, 
      buffer_out_vector_1_55_port, buffer_out_vector_1_54_port, 
      buffer_out_vector_1_53_port, buffer_out_vector_1_52_port, 
      buffer_out_vector_1_51_port, buffer_out_vector_1_50_port, 
      buffer_out_vector_1_49_port, buffer_out_vector_1_48_port, 
      buffer_out_vector_1_47_port, buffer_out_vector_1_46_port, 
      buffer_out_vector_1_45_port, buffer_out_vector_1_44_port, 
      buffer_out_vector_1_43_port, buffer_out_vector_1_42_port, 
      buffer_out_vector_1_41_port, buffer_out_vector_1_40_port, 
      buffer_out_vector_1_39_port, buffer_out_vector_1_38_port, 
      buffer_out_vector_1_37_port, buffer_out_vector_1_36_port, 
      buffer_out_vector_1_35_port, buffer_out_vector_1_34_port, 
      buffer_out_vector_1_33_port, buffer_out_vector_1_32_port, 
      buffer_out_vector_1_31_port, buffer_out_vector_1_30_port, 
      buffer_out_vector_1_29_port, buffer_out_vector_1_28_port, 
      buffer_out_vector_1_27_port, buffer_out_vector_1_26_port, 
      buffer_out_vector_1_25_port, buffer_out_vector_1_24_port, 
      buffer_out_vector_1_23_port, buffer_out_vector_1_22_port, 
      buffer_out_vector_1_21_port, buffer_out_vector_1_20_port, 
      buffer_out_vector_1_19_port, buffer_out_vector_1_18_port, 
      buffer_out_vector_1_17_port, buffer_out_vector_1_16_port, 
      buffer_out_vector_1_15_port, buffer_out_vector_1_14_port, 
      buffer_out_vector_1_13_port, buffer_out_vector_1_12_port, 
      buffer_out_vector_1_11_port, buffer_out_vector_1_10_port, 
      buffer_out_vector_0_63_port, buffer_out_vector_0_62_port, 
      buffer_out_vector_0_61_port, buffer_out_vector_0_60_port, 
      buffer_out_vector_0_59_port, buffer_out_vector_0_58_port, 
      buffer_out_vector_0_57_port, buffer_out_vector_0_56_port, 
      buffer_out_vector_0_55_port, buffer_out_vector_0_54_port, 
      buffer_out_vector_0_53_port, buffer_out_vector_0_52_port, 
      buffer_out_vector_0_51_port, buffer_out_vector_0_50_port, 
      buffer_out_vector_0_49_port, buffer_out_vector_0_48_port, 
      buffer_out_vector_0_47_port, buffer_out_vector_0_46_port, 
      buffer_out_vector_0_45_port, buffer_out_vector_0_44_port, 
      buffer_out_vector_0_43_port, buffer_out_vector_0_42_port, 
      buffer_out_vector_0_41_port, buffer_out_vector_0_40_port, 
      buffer_out_vector_0_39_port, buffer_out_vector_0_38_port, 
      buffer_out_vector_0_37_port, buffer_out_vector_0_36_port, 
      buffer_out_vector_0_35_port, buffer_out_vector_0_34_port, 
      buffer_out_vector_0_33_port, buffer_out_vector_0_32_port, 
      buffer_out_vector_0_31_port, buffer_out_vector_0_30_port, 
      buffer_out_vector_0_29_port, buffer_out_vector_0_28_port, 
      buffer_out_vector_0_27_port, buffer_out_vector_0_26_port, 
      buffer_out_vector_0_25_port, buffer_out_vector_0_24_port, 
      buffer_out_vector_0_23_port, buffer_out_vector_0_22_port, 
      buffer_out_vector_0_21_port, buffer_out_vector_0_20_port, 
      buffer_out_vector_0_19_port, buffer_out_vector_0_18_port, 
      buffer_out_vector_0_17_port, buffer_out_vector_0_16_port, 
      buffer_out_vector_0_15_port, buffer_out_vector_0_14_port, 
      buffer_out_vector_0_13_port, buffer_out_vector_0_12_port, 
      buffer_out_vector_0_11_port, buffer_out_vector_0_10_port, n1, n2, n3, n4,
      n5, n6, n7, n8 : std_logic;

begin
   header <= ( header_1_PACKET_LENGTH_3_port, header_1_PACKET_LENGTH_2_port, 
      header_1_PACKET_LENGTH_1_port, header_1_PACKET_LENGTH_0_port, 
      header_1_X_DEST_1_port, header_1_X_DEST_0_port, header_1_Y_DEST_1_port, 
      header_1_Y_DEST_0_port, header_1_Z_DEST_1_port, header_1_Z_DEST_0_port, 
      header_0_PACKET_LENGTH_3_port, header_0_PACKET_LENGTH_2_port, 
      header_0_PACKET_LENGTH_1_port, header_0_PACKET_LENGTH_0_port, 
      header_0_X_DEST_1_port, header_0_X_DEST_0_port, header_0_Y_DEST_1_port, 
      header_0_Y_DEST_0_port, header_0_Z_DEST_1_port, header_0_Z_DEST_0_port );
   
   U2 : AO22x1_ASAP7_75t_R port map( A1 => n3, A2 => 
                           buffer_out_vector_1_30_port, B1 => 
                           buffer_out_vector_0_30_port, B2 => n4, Y => 
                           data_transfer(30));
   U3 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_31_port, A2 => 
                           n3, B1 => buffer_out_vector_0_31_port, B2 => n4, Y 
                           => data_transfer(31));
   U4 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_32_port, A2 => 
                           n3, B1 => buffer_out_vector_0_32_port, B2 => n4, Y 
                           => data_transfer(32));
   U5 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_33_port, A2 => 
                           n3, B1 => buffer_out_vector_0_33_port, B2 => n4, Y 
                           => data_transfer(33));
   U6 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_34_port, A2 => 
                           n3, B1 => buffer_out_vector_0_34_port, B2 => n4, Y 
                           => data_transfer(34));
   U7 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_35_port, A2 => 
                           n3, B1 => buffer_out_vector_0_35_port, B2 => n7, Y 
                           => data_transfer(35));
   U8 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_36_port, A2 => 
                           n3, B1 => buffer_out_vector_0_36_port, B2 => n6, Y 
                           => data_transfer(36));
   U9 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_37_port, A2 => 
                           n3, B1 => buffer_out_vector_0_37_port, B2 => n7, Y 
                           => data_transfer(37));
   U10 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_38_port, A2 => 
                           n3, B1 => buffer_out_vector_0_38_port, B2 => n5, Y 
                           => data_transfer(38));
   U11 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_39_port, A2 => 
                           n3, B1 => buffer_out_vector_0_39_port, B2 => n7, Y 
                           => data_transfer(39));
   U12 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_40_port, A2 => 
                           n3, B1 => buffer_out_vector_0_40_port, B2 => n6, Y 
                           => data_transfer(40));
   U13 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_41_port, A2 => 
                           n3, B1 => buffer_out_vector_0_41_port, B2 => n5, Y 
                           => data_transfer(41));
   U14 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_42_port, A2 => 
                           n3, B1 => buffer_out_vector_0_42_port, B2 => n5, Y 
                           => data_transfer(42));
   U15 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_43_port, A2 => 
                           n3, B1 => buffer_out_vector_0_43_port, B2 => n5, Y 
                           => data_transfer(43));
   U16 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_44_port, A2 => 
                           n3, B1 => buffer_out_vector_0_44_port, B2 => n7, Y 
                           => data_transfer(44));
   U17 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_45_port, A2 => 
                           n3, B1 => buffer_out_vector_0_45_port, B2 => n5, Y 
                           => data_transfer(45));
   U18 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_46_port, A2 => 
                           n3, B1 => buffer_out_vector_0_46_port, B2 => n6, Y 
                           => data_transfer(46));
   U19 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_47_port, A2 => 
                           n3, B1 => buffer_out_vector_0_47_port, B2 => n7, Y 
                           => data_transfer(47));
   U20 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_48_port, A2 => 
                           n3, B1 => buffer_out_vector_0_48_port, B2 => n6, Y 
                           => data_transfer(48));
   U21 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_49_port, A2 => 
                           n3, B1 => buffer_out_vector_0_49_port, B2 => n7, Y 
                           => data_transfer(49));
   U22 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_50_port, A2 => 
                           n3, B1 => buffer_out_vector_0_50_port, B2 => n5, Y 
                           => data_transfer(50));
   U23 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_51_port, A2 => 
                           n2, B1 => buffer_out_vector_0_51_port, B2 => n5, Y 
                           => data_transfer(51));
   U24 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_52_port, A2 => 
                           n2, B1 => buffer_out_vector_0_52_port, B2 => n7, Y 
                           => data_transfer(52));
   U25 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_53_port, A2 => 
                           n2, B1 => buffer_out_vector_0_53_port, B2 => n6, Y 
                           => data_transfer(53));
   U26 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_54_port, A2 => 
                           n2, B1 => buffer_out_vector_0_54_port, B2 => n6, Y 
                           => data_transfer(54));
   U27 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_55_port, A2 => 
                           n2, B1 => buffer_out_vector_0_55_port, B2 => n7, Y 
                           => data_transfer(55));
   U28 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_56_port, A2 => 
                           n2, B1 => buffer_out_vector_0_56_port, B2 => n6, Y 
                           => data_transfer(56));
   U29 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_57_port, A2 => 
                           n2, B1 => buffer_out_vector_0_57_port, B2 => n6, Y 
                           => data_transfer(57));
   U30 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_58_port, A2 => 
                           n2, B1 => buffer_out_vector_0_58_port, B2 => n5, Y 
                           => data_transfer(58));
   U31 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_59_port, A2 => 
                           n2, B1 => buffer_out_vector_0_59_port, B2 => n5, Y 
                           => data_transfer(59));
   U32 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_60_port, A2 => 
                           n2, B1 => buffer_out_vector_0_60_port, B2 => n5, Y 
                           => data_transfer(60));
   U33 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_61_port, A2 => 
                           n2, B1 => buffer_out_vector_0_61_port, B2 => n5, Y 
                           => data_transfer(61));
   U34 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_62_port, A2 => 
                           n2, B1 => buffer_out_vector_0_62_port, B2 => n5, Y 
                           => data_transfer(62));
   U35 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_63_port, A2 => 
                           n2, B1 => buffer_out_vector_0_63_port, B2 => n5, Y 
                           => data_transfer(63));
   U36 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_0_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_0_port, B2 => n5
                           , Y => data_transfer(0));
   U37 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_1_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_1_port, B2 => n5
                           , Y => data_transfer(1));
   U38 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_2_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_2_port, B2 => n5
                           , Y => data_transfer(2));
   U39 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_3_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_3_port, B2 => n6
                           , Y => data_transfer(3));
   U40 : AO22x1_ASAP7_75t_R port map( A1 => header_1_X_DEST_0_port, A2 => n2, 
                           B1 => header_0_X_DEST_0_port, B2 => n6, Y => 
                           data_transfer(4));
   U41 : AO22x1_ASAP7_75t_R port map( A1 => header_1_X_DEST_1_port, A2 => n2, 
                           B1 => header_0_X_DEST_1_port, B2 => n6, Y => 
                           data_transfer(5));
   U42 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Y_DEST_0_port, A2 => n2, 
                           B1 => header_0_Y_DEST_0_port, B2 => n6, Y => 
                           data_transfer(6));
   U43 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Y_DEST_1_port, A2 => n2, 
                           B1 => header_0_Y_DEST_1_port, B2 => n6, Y => 
                           data_transfer(7));
   U44 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Z_DEST_0_port, A2 => n2, 
                           B1 => header_0_Z_DEST_0_port, B2 => n6, Y => 
                           data_transfer(8));
   U45 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Z_DEST_1_port, A2 => n2, 
                           B1 => header_0_Z_DEST_1_port, B2 => n6, Y => 
                           data_transfer(9));
   U46 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_10_port, A2 => 
                           n2, B1 => buffer_out_vector_0_10_port, B2 => n6, Y 
                           => data_transfer(10));
   U47 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_11_port, A2 => 
                           n2, B1 => buffer_out_vector_0_11_port, B2 => n7, Y 
                           => data_transfer(11));
   U48 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_12_port, A2 => 
                           n2, B1 => buffer_out_vector_0_12_port, B2 => n7, Y 
                           => data_transfer(12));
   U49 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_13_port, A2 => 
                           n2, B1 => buffer_out_vector_0_13_port, B2 => n7, Y 
                           => data_transfer(13));
   U50 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_14_port, A2 => 
                           n2, B1 => buffer_out_vector_0_14_port, B2 => n7, Y 
                           => data_transfer(14));
   U51 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_15_port, A2 => 
                           n2, B1 => buffer_out_vector_0_15_port, B2 => n7, Y 
                           => data_transfer(15));
   U52 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_16_port, A2 => 
                           n2, B1 => buffer_out_vector_0_16_port, B2 => n7, Y 
                           => data_transfer(16));
   U53 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_17_port, A2 => 
                           n2, B1 => buffer_out_vector_0_17_port, B2 => n7, Y 
                           => data_transfer(17));
   U54 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_18_port, A2 => 
                           n2, B1 => buffer_out_vector_0_18_port, B2 => n7, Y 
                           => data_transfer(18));
   U55 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_19_port, A2 => 
                           n2, B1 => buffer_out_vector_0_19_port, B2 => n6, Y 
                           => data_transfer(19));
   U56 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_20_port, A2 => 
                           n2, B1 => buffer_out_vector_0_20_port, B2 => n7, Y 
                           => data_transfer(20));
   U57 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_21_port, A2 => 
                           n2, B1 => buffer_out_vector_0_21_port, B2 => n5, Y 
                           => data_transfer(21));
   U58 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_22_port, A2 => 
                           n2, B1 => buffer_out_vector_0_22_port, B2 => n6, Y 
                           => data_transfer(22));
   U59 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_23_port, A2 => 
                           n2, B1 => buffer_out_vector_0_23_port, B2 => n7, Y 
                           => data_transfer(23));
   U60 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_24_port, A2 => 
                           n2, B1 => buffer_out_vector_0_24_port, B2 => n5, Y 
                           => data_transfer(24));
   U61 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_25_port, A2 => 
                           n2, B1 => buffer_out_vector_0_25_port, B2 => n6, Y 
                           => data_transfer(25));
   U62 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_26_port, A2 => 
                           n2, B1 => buffer_out_vector_0_26_port, B2 => n7, Y 
                           => data_transfer(26));
   U63 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_27_port, A2 => 
                           n2, B1 => buffer_out_vector_0_27_port, B2 => n5, Y 
                           => data_transfer(27));
   U64 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_28_port, A2 => 
                           n2, B1 => buffer_out_vector_0_28_port, B2 => n6, Y 
                           => data_transfer(28));
   U65 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_29_port, A2 => 
                           n2, B1 => buffer_out_vector_0_29_port, B2 => n5, Y 
                           => data_transfer(29));
   fifo_i_0 : fifo_buff_depth2_4 port map( data_in(63) => data_rx(63), 
                           data_in(62) => data_rx(62), data_in(61) => 
                           data_rx(61), data_in(60) => data_rx(60), data_in(59)
                           => data_rx(59), data_in(58) => data_rx(58), 
                           data_in(57) => data_rx(57), data_in(56) => 
                           data_rx(56), data_in(55) => data_rx(55), data_in(54)
                           => data_rx(54), data_in(53) => data_rx(53), 
                           data_in(52) => data_rx(52), data_in(51) => 
                           data_rx(51), data_in(50) => data_rx(50), data_in(49)
                           => data_rx(49), data_in(48) => data_rx(48), 
                           data_in(47) => data_rx(47), data_in(46) => 
                           data_rx(46), data_in(45) => data_rx(45), data_in(44)
                           => data_rx(44), data_in(43) => data_rx(43), 
                           data_in(42) => data_rx(42), data_in(41) => 
                           data_rx(41), data_in(40) => data_rx(40), data_in(39)
                           => data_rx(39), data_in(38) => data_rx(38), 
                           data_in(37) => data_rx(37), data_in(36) => 
                           data_rx(36), data_in(35) => data_rx(35), data_in(34)
                           => data_rx(34), data_in(33) => data_rx(33), 
                           data_in(32) => data_rx(32), data_in(31) => 
                           data_rx(31), data_in(30) => data_rx(30), data_in(29)
                           => data_rx(29), data_in(28) => data_rx(28), 
                           data_in(27) => data_rx(27), data_in(26) => 
                           data_rx(26), data_in(25) => data_rx(25), data_in(24)
                           => data_rx(24), data_in(23) => data_rx(23), 
                           data_in(22) => data_rx(22), data_in(21) => 
                           data_rx(21), data_in(20) => data_rx(20), data_in(19)
                           => data_rx(19), data_in(18) => data_rx(18), 
                           data_in(17) => data_rx(17), data_in(16) => 
                           data_rx(16), data_in(15) => data_rx(15), data_in(14)
                           => data_rx(14), data_in(13) => data_rx(13), 
                           data_in(12) => data_rx(12), data_in(11) => 
                           data_rx(11), data_in(10) => data_rx(10), data_in(9) 
                           => data_rx(9), data_in(8) => data_rx(8), data_in(7) 
                           => data_rx(7), data_in(6) => data_rx(6), data_in(5) 
                           => data_rx(5), data_in(4) => data_rx(4), data_in(3) 
                           => data_rx(3), data_in(2) => data_rx(2), data_in(1) 
                           => data_rx(1), data_in(0) => data_rx(0), write_en =>
                           vc_write_rx(0), read_en => vc_transfer(0), clk => 
                           clk, rst => n8, data_out(63) => 
                           buffer_out_vector_0_63_port, data_out(62) => 
                           buffer_out_vector_0_62_port, data_out(61) => 
                           buffer_out_vector_0_61_port, data_out(60) => 
                           buffer_out_vector_0_60_port, data_out(59) => 
                           buffer_out_vector_0_59_port, data_out(58) => 
                           buffer_out_vector_0_58_port, data_out(57) => 
                           buffer_out_vector_0_57_port, data_out(56) => 
                           buffer_out_vector_0_56_port, data_out(55) => 
                           buffer_out_vector_0_55_port, data_out(54) => 
                           buffer_out_vector_0_54_port, data_out(53) => 
                           buffer_out_vector_0_53_port, data_out(52) => 
                           buffer_out_vector_0_52_port, data_out(51) => 
                           buffer_out_vector_0_51_port, data_out(50) => 
                           buffer_out_vector_0_50_port, data_out(49) => 
                           buffer_out_vector_0_49_port, data_out(48) => 
                           buffer_out_vector_0_48_port, data_out(47) => 
                           buffer_out_vector_0_47_port, data_out(46) => 
                           buffer_out_vector_0_46_port, data_out(45) => 
                           buffer_out_vector_0_45_port, data_out(44) => 
                           buffer_out_vector_0_44_port, data_out(43) => 
                           buffer_out_vector_0_43_port, data_out(42) => 
                           buffer_out_vector_0_42_port, data_out(41) => 
                           buffer_out_vector_0_41_port, data_out(40) => 
                           buffer_out_vector_0_40_port, data_out(39) => 
                           buffer_out_vector_0_39_port, data_out(38) => 
                           buffer_out_vector_0_38_port, data_out(37) => 
                           buffer_out_vector_0_37_port, data_out(36) => 
                           buffer_out_vector_0_36_port, data_out(35) => 
                           buffer_out_vector_0_35_port, data_out(34) => 
                           buffer_out_vector_0_34_port, data_out(33) => 
                           buffer_out_vector_0_33_port, data_out(32) => 
                           buffer_out_vector_0_32_port, data_out(31) => 
                           buffer_out_vector_0_31_port, data_out(30) => 
                           buffer_out_vector_0_30_port, data_out(29) => 
                           buffer_out_vector_0_29_port, data_out(28) => 
                           buffer_out_vector_0_28_port, data_out(27) => 
                           buffer_out_vector_0_27_port, data_out(26) => 
                           buffer_out_vector_0_26_port, data_out(25) => 
                           buffer_out_vector_0_25_port, data_out(24) => 
                           buffer_out_vector_0_24_port, data_out(23) => 
                           buffer_out_vector_0_23_port, data_out(22) => 
                           buffer_out_vector_0_22_port, data_out(21) => 
                           buffer_out_vector_0_21_port, data_out(20) => 
                           buffer_out_vector_0_20_port, data_out(19) => 
                           buffer_out_vector_0_19_port, data_out(18) => 
                           buffer_out_vector_0_18_port, data_out(17) => 
                           buffer_out_vector_0_17_port, data_out(16) => 
                           buffer_out_vector_0_16_port, data_out(15) => 
                           buffer_out_vector_0_15_port, data_out(14) => 
                           buffer_out_vector_0_14_port, data_out(13) => 
                           buffer_out_vector_0_13_port, data_out(12) => 
                           buffer_out_vector_0_12_port, data_out(11) => 
                           buffer_out_vector_0_11_port, data_out(10) => 
                           buffer_out_vector_0_10_port, data_out(9) => 
                           header_0_Z_DEST_1_port, data_out(8) => 
                           header_0_Z_DEST_0_port, data_out(7) => 
                           header_0_Y_DEST_1_port, data_out(6) => 
                           header_0_Y_DEST_0_port, data_out(5) => 
                           header_0_X_DEST_1_port, data_out(4) => 
                           header_0_X_DEST_0_port, data_out(3) => 
                           header_0_PACKET_LENGTH_3_port, data_out(2) => 
                           header_0_PACKET_LENGTH_2_port, data_out(1) => 
                           header_0_PACKET_LENGTH_1_port, data_out(0) => 
                           header_0_PACKET_LENGTH_0_port, valid_data => 
                           valid_data_vc(0));
   fifo_i_1 : fifo_buff_depth2_3 port map( data_in(63) => data_rx(63), 
                           data_in(62) => data_rx(62), data_in(61) => 
                           data_rx(61), data_in(60) => data_rx(60), data_in(59)
                           => data_rx(59), data_in(58) => data_rx(58), 
                           data_in(57) => data_rx(57), data_in(56) => 
                           data_rx(56), data_in(55) => data_rx(55), data_in(54)
                           => data_rx(54), data_in(53) => data_rx(53), 
                           data_in(52) => data_rx(52), data_in(51) => 
                           data_rx(51), data_in(50) => data_rx(50), data_in(49)
                           => data_rx(49), data_in(48) => data_rx(48), 
                           data_in(47) => data_rx(47), data_in(46) => 
                           data_rx(46), data_in(45) => data_rx(45), data_in(44)
                           => data_rx(44), data_in(43) => data_rx(43), 
                           data_in(42) => data_rx(42), data_in(41) => 
                           data_rx(41), data_in(40) => data_rx(40), data_in(39)
                           => data_rx(39), data_in(38) => data_rx(38), 
                           data_in(37) => data_rx(37), data_in(36) => 
                           data_rx(36), data_in(35) => data_rx(35), data_in(34)
                           => data_rx(34), data_in(33) => data_rx(33), 
                           data_in(32) => data_rx(32), data_in(31) => 
                           data_rx(31), data_in(30) => data_rx(30), data_in(29)
                           => data_rx(29), data_in(28) => data_rx(28), 
                           data_in(27) => data_rx(27), data_in(26) => 
                           data_rx(26), data_in(25) => data_rx(25), data_in(24)
                           => data_rx(24), data_in(23) => data_rx(23), 
                           data_in(22) => data_rx(22), data_in(21) => 
                           data_rx(21), data_in(20) => data_rx(20), data_in(19)
                           => data_rx(19), data_in(18) => data_rx(18), 
                           data_in(17) => data_rx(17), data_in(16) => 
                           data_rx(16), data_in(15) => data_rx(15), data_in(14)
                           => data_rx(14), data_in(13) => data_rx(13), 
                           data_in(12) => data_rx(12), data_in(11) => 
                           data_rx(11), data_in(10) => data_rx(10), data_in(9) 
                           => data_rx(9), data_in(8) => data_rx(8), data_in(7) 
                           => data_rx(7), data_in(6) => data_rx(6), data_in(5) 
                           => data_rx(5), data_in(4) => data_rx(4), data_in(3) 
                           => data_rx(3), data_in(2) => data_rx(2), data_in(1) 
                           => data_rx(1), data_in(0) => data_rx(0), write_en =>
                           vc_write_rx(1), read_en => n2, clk => clk, rst => n8
                           , data_out(63) => buffer_out_vector_1_63_port, 
                           data_out(62) => buffer_out_vector_1_62_port, 
                           data_out(61) => buffer_out_vector_1_61_port, 
                           data_out(60) => buffer_out_vector_1_60_port, 
                           data_out(59) => buffer_out_vector_1_59_port, 
                           data_out(58) => buffer_out_vector_1_58_port, 
                           data_out(57) => buffer_out_vector_1_57_port, 
                           data_out(56) => buffer_out_vector_1_56_port, 
                           data_out(55) => buffer_out_vector_1_55_port, 
                           data_out(54) => buffer_out_vector_1_54_port, 
                           data_out(53) => buffer_out_vector_1_53_port, 
                           data_out(52) => buffer_out_vector_1_52_port, 
                           data_out(51) => buffer_out_vector_1_51_port, 
                           data_out(50) => buffer_out_vector_1_50_port, 
                           data_out(49) => buffer_out_vector_1_49_port, 
                           data_out(48) => buffer_out_vector_1_48_port, 
                           data_out(47) => buffer_out_vector_1_47_port, 
                           data_out(46) => buffer_out_vector_1_46_port, 
                           data_out(45) => buffer_out_vector_1_45_port, 
                           data_out(44) => buffer_out_vector_1_44_port, 
                           data_out(43) => buffer_out_vector_1_43_port, 
                           data_out(42) => buffer_out_vector_1_42_port, 
                           data_out(41) => buffer_out_vector_1_41_port, 
                           data_out(40) => buffer_out_vector_1_40_port, 
                           data_out(39) => buffer_out_vector_1_39_port, 
                           data_out(38) => buffer_out_vector_1_38_port, 
                           data_out(37) => buffer_out_vector_1_37_port, 
                           data_out(36) => buffer_out_vector_1_36_port, 
                           data_out(35) => buffer_out_vector_1_35_port, 
                           data_out(34) => buffer_out_vector_1_34_port, 
                           data_out(33) => buffer_out_vector_1_33_port, 
                           data_out(32) => buffer_out_vector_1_32_port, 
                           data_out(31) => buffer_out_vector_1_31_port, 
                           data_out(30) => buffer_out_vector_1_30_port, 
                           data_out(29) => buffer_out_vector_1_29_port, 
                           data_out(28) => buffer_out_vector_1_28_port, 
                           data_out(27) => buffer_out_vector_1_27_port, 
                           data_out(26) => buffer_out_vector_1_26_port, 
                           data_out(25) => buffer_out_vector_1_25_port, 
                           data_out(24) => buffer_out_vector_1_24_port, 
                           data_out(23) => buffer_out_vector_1_23_port, 
                           data_out(22) => buffer_out_vector_1_22_port, 
                           data_out(21) => buffer_out_vector_1_21_port, 
                           data_out(20) => buffer_out_vector_1_20_port, 
                           data_out(19) => buffer_out_vector_1_19_port, 
                           data_out(18) => buffer_out_vector_1_18_port, 
                           data_out(17) => buffer_out_vector_1_17_port, 
                           data_out(16) => buffer_out_vector_1_16_port, 
                           data_out(15) => buffer_out_vector_1_15_port, 
                           data_out(14) => buffer_out_vector_1_14_port, 
                           data_out(13) => buffer_out_vector_1_13_port, 
                           data_out(12) => buffer_out_vector_1_12_port, 
                           data_out(11) => buffer_out_vector_1_11_port, 
                           data_out(10) => buffer_out_vector_1_10_port, 
                           data_out(9) => header_1_Z_DEST_1_port, data_out(8) 
                           => header_1_Z_DEST_0_port, data_out(7) => 
                           header_1_Y_DEST_1_port, data_out(6) => 
                           header_1_Y_DEST_0_port, data_out(5) => 
                           header_1_X_DEST_1_port, data_out(4) => 
                           header_1_X_DEST_0_port, data_out(3) => 
                           header_1_PACKET_LENGTH_3_port, data_out(2) => 
                           header_1_PACKET_LENGTH_2_port, data_out(1) => 
                           header_1_PACKET_LENGTH_1_port, data_out(0) => 
                           header_1_PACKET_LENGTH_0_port, valid_data => 
                           valid_data_vc(1));
   U1 : INVx1_ASAP7_75t_R port map( A => n4, Y => n2);
   U66 : INVx1_ASAP7_75t_R port map( A => n4, Y => n3);
   U67 : INVx1_ASAP7_75t_R port map( A => n1, Y => n4);
   U68 : INVx1_ASAP7_75t_R port map( A => n1, Y => n6);
   U69 : INVx1_ASAP7_75t_R port map( A => n1, Y => n5);
   U70 : INVx1_ASAP7_75t_R port map( A => n1, Y => n7);
   U71 : HB1xp67_ASAP7_75t_R port map( A => vc_transfer(1), Y => n1);
   U72 : HB1xp67_ASAP7_75t_R port map( A => rst, Y => n8);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity vc_input_buffer_2_0000000200000002_1 is

   port( clk, rst : in std_logic;  data_rx : in std_logic_vector (63 downto 0);
         vc_write_rx, vc_transfer : in std_logic_vector (1 downto 0);  
         valid_data_vc : out std_logic_vector (1 downto 0);  data_transfer : 
         out std_logic_vector (63 downto 0);  header : out std_logic_vector (19
         downto 0));

end vc_input_buffer_2_0000000200000002_1;

architecture SYN_rtl of vc_input_buffer_2_0000000200000002_1 is

   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component fifo_buff_depth2_1
      port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, 
            clk, rst : in std_logic;  data_out : out std_logic_vector (63 
            downto 0);  valid_data : out std_logic);
   end component;
   
   component fifo_buff_depth2_2
      port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, 
            clk, rst : in std_logic;  data_out : out std_logic_vector (63 
            downto 0);  valid_data : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal header_1_PACKET_LENGTH_3_port, header_1_PACKET_LENGTH_2_port, 
      header_1_PACKET_LENGTH_1_port, header_1_PACKET_LENGTH_0_port, 
      header_1_X_DEST_1_port, header_1_X_DEST_0_port, header_1_Y_DEST_1_port, 
      header_1_Y_DEST_0_port, header_1_Z_DEST_1_port, header_1_Z_DEST_0_port, 
      header_0_PACKET_LENGTH_3_port, header_0_PACKET_LENGTH_2_port, 
      header_0_PACKET_LENGTH_1_port, header_0_PACKET_LENGTH_0_port, 
      header_0_X_DEST_1_port, header_0_X_DEST_0_port, header_0_Y_DEST_1_port, 
      header_0_Y_DEST_0_port, header_0_Z_DEST_1_port, header_0_Z_DEST_0_port, 
      buffer_out_vector_1_63_port, buffer_out_vector_1_62_port, 
      buffer_out_vector_1_61_port, buffer_out_vector_1_60_port, 
      buffer_out_vector_1_59_port, buffer_out_vector_1_58_port, 
      buffer_out_vector_1_57_port, buffer_out_vector_1_56_port, 
      buffer_out_vector_1_55_port, buffer_out_vector_1_54_port, 
      buffer_out_vector_1_53_port, buffer_out_vector_1_52_port, 
      buffer_out_vector_1_51_port, buffer_out_vector_1_50_port, 
      buffer_out_vector_1_49_port, buffer_out_vector_1_48_port, 
      buffer_out_vector_1_47_port, buffer_out_vector_1_46_port, 
      buffer_out_vector_1_45_port, buffer_out_vector_1_44_port, 
      buffer_out_vector_1_43_port, buffer_out_vector_1_42_port, 
      buffer_out_vector_1_41_port, buffer_out_vector_1_40_port, 
      buffer_out_vector_1_39_port, buffer_out_vector_1_38_port, 
      buffer_out_vector_1_37_port, buffer_out_vector_1_36_port, 
      buffer_out_vector_1_35_port, buffer_out_vector_1_34_port, 
      buffer_out_vector_1_33_port, buffer_out_vector_1_32_port, 
      buffer_out_vector_1_31_port, buffer_out_vector_1_30_port, 
      buffer_out_vector_1_29_port, buffer_out_vector_1_28_port, 
      buffer_out_vector_1_27_port, buffer_out_vector_1_26_port, 
      buffer_out_vector_1_25_port, buffer_out_vector_1_24_port, 
      buffer_out_vector_1_23_port, buffer_out_vector_1_22_port, 
      buffer_out_vector_1_21_port, buffer_out_vector_1_20_port, 
      buffer_out_vector_1_19_port, buffer_out_vector_1_18_port, 
      buffer_out_vector_1_17_port, buffer_out_vector_1_16_port, 
      buffer_out_vector_1_15_port, buffer_out_vector_1_14_port, 
      buffer_out_vector_1_13_port, buffer_out_vector_1_12_port, 
      buffer_out_vector_1_11_port, buffer_out_vector_1_10_port, 
      buffer_out_vector_0_63_port, buffer_out_vector_0_62_port, 
      buffer_out_vector_0_61_port, buffer_out_vector_0_60_port, 
      buffer_out_vector_0_59_port, buffer_out_vector_0_58_port, 
      buffer_out_vector_0_57_port, buffer_out_vector_0_56_port, 
      buffer_out_vector_0_55_port, buffer_out_vector_0_54_port, 
      buffer_out_vector_0_53_port, buffer_out_vector_0_52_port, 
      buffer_out_vector_0_51_port, buffer_out_vector_0_50_port, 
      buffer_out_vector_0_49_port, buffer_out_vector_0_48_port, 
      buffer_out_vector_0_47_port, buffer_out_vector_0_46_port, 
      buffer_out_vector_0_45_port, buffer_out_vector_0_44_port, 
      buffer_out_vector_0_43_port, buffer_out_vector_0_42_port, 
      buffer_out_vector_0_41_port, buffer_out_vector_0_40_port, 
      buffer_out_vector_0_39_port, buffer_out_vector_0_38_port, 
      buffer_out_vector_0_37_port, buffer_out_vector_0_36_port, 
      buffer_out_vector_0_35_port, buffer_out_vector_0_34_port, 
      buffer_out_vector_0_33_port, buffer_out_vector_0_32_port, 
      buffer_out_vector_0_31_port, buffer_out_vector_0_30_port, 
      buffer_out_vector_0_29_port, buffer_out_vector_0_28_port, 
      buffer_out_vector_0_27_port, buffer_out_vector_0_26_port, 
      buffer_out_vector_0_25_port, buffer_out_vector_0_24_port, 
      buffer_out_vector_0_23_port, buffer_out_vector_0_22_port, 
      buffer_out_vector_0_21_port, buffer_out_vector_0_20_port, 
      buffer_out_vector_0_19_port, buffer_out_vector_0_18_port, 
      buffer_out_vector_0_17_port, buffer_out_vector_0_16_port, 
      buffer_out_vector_0_15_port, buffer_out_vector_0_14_port, 
      buffer_out_vector_0_13_port, buffer_out_vector_0_12_port, 
      buffer_out_vector_0_11_port, buffer_out_vector_0_10_port, n1, n2, n3, n4,
      n5, n6, n7 : std_logic;

begin
   header <= ( header_1_PACKET_LENGTH_3_port, header_1_PACKET_LENGTH_2_port, 
      header_1_PACKET_LENGTH_1_port, header_1_PACKET_LENGTH_0_port, 
      header_1_X_DEST_1_port, header_1_X_DEST_0_port, header_1_Y_DEST_1_port, 
      header_1_Y_DEST_0_port, header_1_Z_DEST_1_port, header_1_Z_DEST_0_port, 
      header_0_PACKET_LENGTH_3_port, header_0_PACKET_LENGTH_2_port, 
      header_0_PACKET_LENGTH_1_port, header_0_PACKET_LENGTH_0_port, 
      header_0_X_DEST_1_port, header_0_X_DEST_0_port, header_0_Y_DEST_1_port, 
      header_0_Y_DEST_0_port, header_0_Z_DEST_1_port, header_0_Z_DEST_0_port );
   
   U2 : AO22x1_ASAP7_75t_R port map( A1 => n3, A2 => 
                           buffer_out_vector_1_30_port, B1 => 
                           buffer_out_vector_0_30_port, B2 => n4, Y => 
                           data_transfer(30));
   U3 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_31_port, A2 => 
                           n3, B1 => buffer_out_vector_0_31_port, B2 => n4, Y 
                           => data_transfer(31));
   U4 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_32_port, A2 => 
                           n3, B1 => buffer_out_vector_0_32_port, B2 => n4, Y 
                           => data_transfer(32));
   U5 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_33_port, A2 => 
                           n3, B1 => buffer_out_vector_0_33_port, B2 => n4, Y 
                           => data_transfer(33));
   U6 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_34_port, A2 => 
                           n3, B1 => buffer_out_vector_0_34_port, B2 => n4, Y 
                           => data_transfer(34));
   U7 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_35_port, A2 => 
                           n3, B1 => buffer_out_vector_0_35_port, B2 => n6, Y 
                           => data_transfer(35));
   U8 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_36_port, A2 => 
                           n3, B1 => buffer_out_vector_0_36_port, B2 => n6, Y 
                           => data_transfer(36));
   U9 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_37_port, A2 => 
                           n3, B1 => buffer_out_vector_0_37_port, B2 => n5, Y 
                           => data_transfer(37));
   U10 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_38_port, A2 => 
                           n3, B1 => buffer_out_vector_0_38_port, B2 => n5, Y 
                           => data_transfer(38));
   U11 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_39_port, A2 => 
                           n3, B1 => buffer_out_vector_0_39_port, B2 => n5, Y 
                           => data_transfer(39));
   U12 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_40_port, A2 => 
                           n3, B1 => buffer_out_vector_0_40_port, B2 => n6, Y 
                           => data_transfer(40));
   U13 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_41_port, A2 => 
                           n3, B1 => buffer_out_vector_0_41_port, B2 => n5, Y 
                           => data_transfer(41));
   U14 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_42_port, A2 => 
                           n3, B1 => buffer_out_vector_0_42_port, B2 => n5, Y 
                           => data_transfer(42));
   U15 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_43_port, A2 => 
                           n3, B1 => buffer_out_vector_0_43_port, B2 => n5, Y 
                           => data_transfer(43));
   U16 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_44_port, A2 => 
                           n3, B1 => buffer_out_vector_0_44_port, B2 => n6, Y 
                           => data_transfer(44));
   U17 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_45_port, A2 => 
                           n3, B1 => buffer_out_vector_0_45_port, B2 => n5, Y 
                           => data_transfer(45));
   U18 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_46_port, A2 => 
                           n3, B1 => buffer_out_vector_0_46_port, B2 => n6, Y 
                           => data_transfer(46));
   U19 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_47_port, A2 => 
                           n3, B1 => buffer_out_vector_0_47_port, B2 => n6, Y 
                           => data_transfer(47));
   U20 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_48_port, A2 => 
                           n3, B1 => buffer_out_vector_0_48_port, B2 => n6, Y 
                           => data_transfer(48));
   U21 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_49_port, A2 => 
                           n3, B1 => buffer_out_vector_0_49_port, B2 => n5, Y 
                           => data_transfer(49));
   U22 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_50_port, A2 => 
                           n3, B1 => buffer_out_vector_0_50_port, B2 => n5, Y 
                           => data_transfer(50));
   U23 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_51_port, A2 => 
                           n2, B1 => buffer_out_vector_0_51_port, B2 => n5, Y 
                           => data_transfer(51));
   U24 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_52_port, A2 => 
                           n2, B1 => buffer_out_vector_0_52_port, B2 => n6, Y 
                           => data_transfer(52));
   U25 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_53_port, A2 => 
                           n2, B1 => buffer_out_vector_0_53_port, B2 => n6, Y 
                           => data_transfer(53));
   U26 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_54_port, A2 => 
                           n2, B1 => buffer_out_vector_0_54_port, B2 => n6, Y 
                           => data_transfer(54));
   U27 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_55_port, A2 => 
                           n2, B1 => buffer_out_vector_0_55_port, B2 => n5, Y 
                           => data_transfer(55));
   U28 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_56_port, A2 => 
                           n2, B1 => buffer_out_vector_0_56_port, B2 => n6, Y 
                           => data_transfer(56));
   U29 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_57_port, A2 => 
                           n2, B1 => buffer_out_vector_0_57_port, B2 => n6, Y 
                           => data_transfer(57));
   U30 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_58_port, A2 => 
                           n2, B1 => buffer_out_vector_0_58_port, B2 => n5, Y 
                           => data_transfer(58));
   U31 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_59_port, A2 => 
                           n2, B1 => buffer_out_vector_0_59_port, B2 => n5, Y 
                           => data_transfer(59));
   U32 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_60_port, A2 => 
                           n2, B1 => buffer_out_vector_0_60_port, B2 => n5, Y 
                           => data_transfer(60));
   U33 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_61_port, A2 => 
                           n2, B1 => buffer_out_vector_0_61_port, B2 => n5, Y 
                           => data_transfer(61));
   U34 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_62_port, A2 => 
                           n2, B1 => buffer_out_vector_0_62_port, B2 => n5, Y 
                           => data_transfer(62));
   U35 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_63_port, A2 => 
                           n2, B1 => buffer_out_vector_0_63_port, B2 => n5, Y 
                           => data_transfer(63));
   U36 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_0_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_0_port, B2 => n5
                           , Y => data_transfer(0));
   U37 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_1_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_1_port, B2 => n5
                           , Y => data_transfer(1));
   U38 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_2_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_2_port, B2 => n5
                           , Y => data_transfer(2));
   U39 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_3_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_3_port, B2 => n6
                           , Y => data_transfer(3));
   U40 : AO22x1_ASAP7_75t_R port map( A1 => header_1_X_DEST_0_port, A2 => n2, 
                           B1 => header_0_X_DEST_0_port, B2 => n6, Y => 
                           data_transfer(4));
   U41 : AO22x1_ASAP7_75t_R port map( A1 => header_1_X_DEST_1_port, A2 => n2, 
                           B1 => header_0_X_DEST_1_port, B2 => n6, Y => 
                           data_transfer(5));
   U42 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Y_DEST_0_port, A2 => n2, 
                           B1 => header_0_Y_DEST_0_port, B2 => n6, Y => 
                           data_transfer(6));
   U43 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Y_DEST_1_port, A2 => n2, 
                           B1 => header_0_Y_DEST_1_port, B2 => n6, Y => 
                           data_transfer(7));
   U44 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Z_DEST_0_port, A2 => n2, 
                           B1 => header_0_Z_DEST_0_port, B2 => n6, Y => 
                           data_transfer(8));
   U45 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Z_DEST_1_port, A2 => n2, 
                           B1 => header_0_Z_DEST_1_port, B2 => n6, Y => 
                           data_transfer(9));
   U46 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_10_port, A2 => 
                           n2, B1 => buffer_out_vector_0_10_port, B2 => n6, Y 
                           => data_transfer(10));
   U47 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_11_port, A2 => 
                           n2, B1 => buffer_out_vector_0_11_port, B2 => n6, Y 
                           => data_transfer(11));
   U48 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_12_port, A2 => 
                           n2, B1 => buffer_out_vector_0_12_port, B2 => n5, Y 
                           => data_transfer(12));
   U49 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_13_port, A2 => 
                           n2, B1 => buffer_out_vector_0_13_port, B2 => n6, Y 
                           => data_transfer(13));
   U50 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_14_port, A2 => 
                           n2, B1 => buffer_out_vector_0_14_port, B2 => n5, Y 
                           => data_transfer(14));
   U51 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_15_port, A2 => 
                           n2, B1 => buffer_out_vector_0_15_port, B2 => n6, Y 
                           => data_transfer(15));
   U52 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_16_port, A2 => 
                           n2, B1 => buffer_out_vector_0_16_port, B2 => n5, Y 
                           => data_transfer(16));
   U53 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_17_port, A2 => 
                           n2, B1 => buffer_out_vector_0_17_port, B2 => n6, Y 
                           => data_transfer(17));
   U54 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_18_port, A2 => 
                           n2, B1 => buffer_out_vector_0_18_port, B2 => n5, Y 
                           => data_transfer(18));
   U55 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_19_port, A2 => 
                           n2, B1 => buffer_out_vector_0_19_port, B2 => n6, Y 
                           => data_transfer(19));
   U56 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_20_port, A2 => 
                           n2, B1 => buffer_out_vector_0_20_port, B2 => n6, Y 
                           => data_transfer(20));
   U57 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_21_port, A2 => 
                           n2, B1 => buffer_out_vector_0_21_port, B2 => n5, Y 
                           => data_transfer(21));
   U58 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_22_port, A2 => 
                           n2, B1 => buffer_out_vector_0_22_port, B2 => n6, Y 
                           => data_transfer(22));
   U59 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_23_port, A2 => 
                           n2, B1 => buffer_out_vector_0_23_port, B2 => n5, Y 
                           => data_transfer(23));
   U60 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_24_port, A2 => 
                           n2, B1 => buffer_out_vector_0_24_port, B2 => n5, Y 
                           => data_transfer(24));
   U61 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_25_port, A2 => 
                           n2, B1 => buffer_out_vector_0_25_port, B2 => n6, Y 
                           => data_transfer(25));
   U62 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_26_port, A2 => 
                           n2, B1 => buffer_out_vector_0_26_port, B2 => n6, Y 
                           => data_transfer(26));
   U63 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_27_port, A2 => 
                           n2, B1 => buffer_out_vector_0_27_port, B2 => n5, Y 
                           => data_transfer(27));
   U64 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_28_port, A2 => 
                           n2, B1 => buffer_out_vector_0_28_port, B2 => n6, Y 
                           => data_transfer(28));
   U65 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_29_port, A2 => 
                           n2, B1 => buffer_out_vector_0_29_port, B2 => n5, Y 
                           => data_transfer(29));
   fifo_i_0 : fifo_buff_depth2_2 port map( data_in(63) => data_rx(63), 
                           data_in(62) => data_rx(62), data_in(61) => 
                           data_rx(61), data_in(60) => data_rx(60), data_in(59)
                           => data_rx(59), data_in(58) => data_rx(58), 
                           data_in(57) => data_rx(57), data_in(56) => 
                           data_rx(56), data_in(55) => data_rx(55), data_in(54)
                           => data_rx(54), data_in(53) => data_rx(53), 
                           data_in(52) => data_rx(52), data_in(51) => 
                           data_rx(51), data_in(50) => data_rx(50), data_in(49)
                           => data_rx(49), data_in(48) => data_rx(48), 
                           data_in(47) => data_rx(47), data_in(46) => 
                           data_rx(46), data_in(45) => data_rx(45), data_in(44)
                           => data_rx(44), data_in(43) => data_rx(43), 
                           data_in(42) => data_rx(42), data_in(41) => 
                           data_rx(41), data_in(40) => data_rx(40), data_in(39)
                           => data_rx(39), data_in(38) => data_rx(38), 
                           data_in(37) => data_rx(37), data_in(36) => 
                           data_rx(36), data_in(35) => data_rx(35), data_in(34)
                           => data_rx(34), data_in(33) => data_rx(33), 
                           data_in(32) => data_rx(32), data_in(31) => 
                           data_rx(31), data_in(30) => data_rx(30), data_in(29)
                           => data_rx(29), data_in(28) => data_rx(28), 
                           data_in(27) => data_rx(27), data_in(26) => 
                           data_rx(26), data_in(25) => data_rx(25), data_in(24)
                           => data_rx(24), data_in(23) => data_rx(23), 
                           data_in(22) => data_rx(22), data_in(21) => 
                           data_rx(21), data_in(20) => data_rx(20), data_in(19)
                           => data_rx(19), data_in(18) => data_rx(18), 
                           data_in(17) => data_rx(17), data_in(16) => 
                           data_rx(16), data_in(15) => data_rx(15), data_in(14)
                           => data_rx(14), data_in(13) => data_rx(13), 
                           data_in(12) => data_rx(12), data_in(11) => 
                           data_rx(11), data_in(10) => data_rx(10), data_in(9) 
                           => data_rx(9), data_in(8) => data_rx(8), data_in(7) 
                           => data_rx(7), data_in(6) => data_rx(6), data_in(5) 
                           => data_rx(5), data_in(4) => data_rx(4), data_in(3) 
                           => data_rx(3), data_in(2) => data_rx(2), data_in(1) 
                           => data_rx(1), data_in(0) => data_rx(0), write_en =>
                           vc_write_rx(0), read_en => vc_transfer(0), clk => 
                           clk, rst => n7, data_out(63) => 
                           buffer_out_vector_0_63_port, data_out(62) => 
                           buffer_out_vector_0_62_port, data_out(61) => 
                           buffer_out_vector_0_61_port, data_out(60) => 
                           buffer_out_vector_0_60_port, data_out(59) => 
                           buffer_out_vector_0_59_port, data_out(58) => 
                           buffer_out_vector_0_58_port, data_out(57) => 
                           buffer_out_vector_0_57_port, data_out(56) => 
                           buffer_out_vector_0_56_port, data_out(55) => 
                           buffer_out_vector_0_55_port, data_out(54) => 
                           buffer_out_vector_0_54_port, data_out(53) => 
                           buffer_out_vector_0_53_port, data_out(52) => 
                           buffer_out_vector_0_52_port, data_out(51) => 
                           buffer_out_vector_0_51_port, data_out(50) => 
                           buffer_out_vector_0_50_port, data_out(49) => 
                           buffer_out_vector_0_49_port, data_out(48) => 
                           buffer_out_vector_0_48_port, data_out(47) => 
                           buffer_out_vector_0_47_port, data_out(46) => 
                           buffer_out_vector_0_46_port, data_out(45) => 
                           buffer_out_vector_0_45_port, data_out(44) => 
                           buffer_out_vector_0_44_port, data_out(43) => 
                           buffer_out_vector_0_43_port, data_out(42) => 
                           buffer_out_vector_0_42_port, data_out(41) => 
                           buffer_out_vector_0_41_port, data_out(40) => 
                           buffer_out_vector_0_40_port, data_out(39) => 
                           buffer_out_vector_0_39_port, data_out(38) => 
                           buffer_out_vector_0_38_port, data_out(37) => 
                           buffer_out_vector_0_37_port, data_out(36) => 
                           buffer_out_vector_0_36_port, data_out(35) => 
                           buffer_out_vector_0_35_port, data_out(34) => 
                           buffer_out_vector_0_34_port, data_out(33) => 
                           buffer_out_vector_0_33_port, data_out(32) => 
                           buffer_out_vector_0_32_port, data_out(31) => 
                           buffer_out_vector_0_31_port, data_out(30) => 
                           buffer_out_vector_0_30_port, data_out(29) => 
                           buffer_out_vector_0_29_port, data_out(28) => 
                           buffer_out_vector_0_28_port, data_out(27) => 
                           buffer_out_vector_0_27_port, data_out(26) => 
                           buffer_out_vector_0_26_port, data_out(25) => 
                           buffer_out_vector_0_25_port, data_out(24) => 
                           buffer_out_vector_0_24_port, data_out(23) => 
                           buffer_out_vector_0_23_port, data_out(22) => 
                           buffer_out_vector_0_22_port, data_out(21) => 
                           buffer_out_vector_0_21_port, data_out(20) => 
                           buffer_out_vector_0_20_port, data_out(19) => 
                           buffer_out_vector_0_19_port, data_out(18) => 
                           buffer_out_vector_0_18_port, data_out(17) => 
                           buffer_out_vector_0_17_port, data_out(16) => 
                           buffer_out_vector_0_16_port, data_out(15) => 
                           buffer_out_vector_0_15_port, data_out(14) => 
                           buffer_out_vector_0_14_port, data_out(13) => 
                           buffer_out_vector_0_13_port, data_out(12) => 
                           buffer_out_vector_0_12_port, data_out(11) => 
                           buffer_out_vector_0_11_port, data_out(10) => 
                           buffer_out_vector_0_10_port, data_out(9) => 
                           header_0_Z_DEST_1_port, data_out(8) => 
                           header_0_Z_DEST_0_port, data_out(7) => 
                           header_0_Y_DEST_1_port, data_out(6) => 
                           header_0_Y_DEST_0_port, data_out(5) => 
                           header_0_X_DEST_1_port, data_out(4) => 
                           header_0_X_DEST_0_port, data_out(3) => 
                           header_0_PACKET_LENGTH_3_port, data_out(2) => 
                           header_0_PACKET_LENGTH_2_port, data_out(1) => 
                           header_0_PACKET_LENGTH_1_port, data_out(0) => 
                           header_0_PACKET_LENGTH_0_port, valid_data => 
                           valid_data_vc(0));
   fifo_i_1 : fifo_buff_depth2_1 port map( data_in(63) => data_rx(63), 
                           data_in(62) => data_rx(62), data_in(61) => 
                           data_rx(61), data_in(60) => data_rx(60), data_in(59)
                           => data_rx(59), data_in(58) => data_rx(58), 
                           data_in(57) => data_rx(57), data_in(56) => 
                           data_rx(56), data_in(55) => data_rx(55), data_in(54)
                           => data_rx(54), data_in(53) => data_rx(53), 
                           data_in(52) => data_rx(52), data_in(51) => 
                           data_rx(51), data_in(50) => data_rx(50), data_in(49)
                           => data_rx(49), data_in(48) => data_rx(48), 
                           data_in(47) => data_rx(47), data_in(46) => 
                           data_rx(46), data_in(45) => data_rx(45), data_in(44)
                           => data_rx(44), data_in(43) => data_rx(43), 
                           data_in(42) => data_rx(42), data_in(41) => 
                           data_rx(41), data_in(40) => data_rx(40), data_in(39)
                           => data_rx(39), data_in(38) => data_rx(38), 
                           data_in(37) => data_rx(37), data_in(36) => 
                           data_rx(36), data_in(35) => data_rx(35), data_in(34)
                           => data_rx(34), data_in(33) => data_rx(33), 
                           data_in(32) => data_rx(32), data_in(31) => 
                           data_rx(31), data_in(30) => data_rx(30), data_in(29)
                           => data_rx(29), data_in(28) => data_rx(28), 
                           data_in(27) => data_rx(27), data_in(26) => 
                           data_rx(26), data_in(25) => data_rx(25), data_in(24)
                           => data_rx(24), data_in(23) => data_rx(23), 
                           data_in(22) => data_rx(22), data_in(21) => 
                           data_rx(21), data_in(20) => data_rx(20), data_in(19)
                           => data_rx(19), data_in(18) => data_rx(18), 
                           data_in(17) => data_rx(17), data_in(16) => 
                           data_rx(16), data_in(15) => data_rx(15), data_in(14)
                           => data_rx(14), data_in(13) => data_rx(13), 
                           data_in(12) => data_rx(12), data_in(11) => 
                           data_rx(11), data_in(10) => data_rx(10), data_in(9) 
                           => data_rx(9), data_in(8) => data_rx(8), data_in(7) 
                           => data_rx(7), data_in(6) => data_rx(6), data_in(5) 
                           => data_rx(5), data_in(4) => data_rx(4), data_in(3) 
                           => data_rx(3), data_in(2) => data_rx(2), data_in(1) 
                           => data_rx(1), data_in(0) => data_rx(0), write_en =>
                           vc_write_rx(1), read_en => n2, clk => clk, rst => n7
                           , data_out(63) => buffer_out_vector_1_63_port, 
                           data_out(62) => buffer_out_vector_1_62_port, 
                           data_out(61) => buffer_out_vector_1_61_port, 
                           data_out(60) => buffer_out_vector_1_60_port, 
                           data_out(59) => buffer_out_vector_1_59_port, 
                           data_out(58) => buffer_out_vector_1_58_port, 
                           data_out(57) => buffer_out_vector_1_57_port, 
                           data_out(56) => buffer_out_vector_1_56_port, 
                           data_out(55) => buffer_out_vector_1_55_port, 
                           data_out(54) => buffer_out_vector_1_54_port, 
                           data_out(53) => buffer_out_vector_1_53_port, 
                           data_out(52) => buffer_out_vector_1_52_port, 
                           data_out(51) => buffer_out_vector_1_51_port, 
                           data_out(50) => buffer_out_vector_1_50_port, 
                           data_out(49) => buffer_out_vector_1_49_port, 
                           data_out(48) => buffer_out_vector_1_48_port, 
                           data_out(47) => buffer_out_vector_1_47_port, 
                           data_out(46) => buffer_out_vector_1_46_port, 
                           data_out(45) => buffer_out_vector_1_45_port, 
                           data_out(44) => buffer_out_vector_1_44_port, 
                           data_out(43) => buffer_out_vector_1_43_port, 
                           data_out(42) => buffer_out_vector_1_42_port, 
                           data_out(41) => buffer_out_vector_1_41_port, 
                           data_out(40) => buffer_out_vector_1_40_port, 
                           data_out(39) => buffer_out_vector_1_39_port, 
                           data_out(38) => buffer_out_vector_1_38_port, 
                           data_out(37) => buffer_out_vector_1_37_port, 
                           data_out(36) => buffer_out_vector_1_36_port, 
                           data_out(35) => buffer_out_vector_1_35_port, 
                           data_out(34) => buffer_out_vector_1_34_port, 
                           data_out(33) => buffer_out_vector_1_33_port, 
                           data_out(32) => buffer_out_vector_1_32_port, 
                           data_out(31) => buffer_out_vector_1_31_port, 
                           data_out(30) => buffer_out_vector_1_30_port, 
                           data_out(29) => buffer_out_vector_1_29_port, 
                           data_out(28) => buffer_out_vector_1_28_port, 
                           data_out(27) => buffer_out_vector_1_27_port, 
                           data_out(26) => buffer_out_vector_1_26_port, 
                           data_out(25) => buffer_out_vector_1_25_port, 
                           data_out(24) => buffer_out_vector_1_24_port, 
                           data_out(23) => buffer_out_vector_1_23_port, 
                           data_out(22) => buffer_out_vector_1_22_port, 
                           data_out(21) => buffer_out_vector_1_21_port, 
                           data_out(20) => buffer_out_vector_1_20_port, 
                           data_out(19) => buffer_out_vector_1_19_port, 
                           data_out(18) => buffer_out_vector_1_18_port, 
                           data_out(17) => buffer_out_vector_1_17_port, 
                           data_out(16) => buffer_out_vector_1_16_port, 
                           data_out(15) => buffer_out_vector_1_15_port, 
                           data_out(14) => buffer_out_vector_1_14_port, 
                           data_out(13) => buffer_out_vector_1_13_port, 
                           data_out(12) => buffer_out_vector_1_12_port, 
                           data_out(11) => buffer_out_vector_1_11_port, 
                           data_out(10) => buffer_out_vector_1_10_port, 
                           data_out(9) => header_1_Z_DEST_1_port, data_out(8) 
                           => header_1_Z_DEST_0_port, data_out(7) => 
                           header_1_Y_DEST_1_port, data_out(6) => 
                           header_1_Y_DEST_0_port, data_out(5) => 
                           header_1_X_DEST_1_port, data_out(4) => 
                           header_1_X_DEST_0_port, data_out(3) => 
                           header_1_PACKET_LENGTH_3_port, data_out(2) => 
                           header_1_PACKET_LENGTH_2_port, data_out(1) => 
                           header_1_PACKET_LENGTH_1_port, data_out(0) => 
                           header_1_PACKET_LENGTH_0_port, valid_data => 
                           valid_data_vc(1));
   U1 : INVx1_ASAP7_75t_R port map( A => n4, Y => n2);
   U66 : INVx1_ASAP7_75t_R port map( A => n4, Y => n3);
   U67 : INVx1_ASAP7_75t_R port map( A => n1, Y => n4);
   U68 : INVx1_ASAP7_75t_R port map( A => n1, Y => n6);
   U69 : INVx1_ASAP7_75t_R port map( A => n1, Y => n5);
   U70 : HB1xp67_ASAP7_75t_R port map( A => vc_transfer(1), Y => n1);
   U71 : HB1xp67_ASAP7_75t_R port map( A => rst, Y => n7);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity dxyu_routing_Xis1_Yis1_Zis1_0 is

   port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;  
         routing : out std_logic_vector (6 downto 0));

end dxyu_routing_Xis1_Yis1_Zis1_0;

architecture SYN_rtl of dxyu_routing_Xis1_Yis1_Zis1_0 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n20, n21, n22, n23, n24, n1, n2, n3, n4, n5, n6, n7 : std_logic;

begin
   
   U8 : NAND2xp5_ASAP7_75t_R port map( A => enable, B => n6, Y => n23);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => n3, B => n2, Y => n22);
   U19 : AND2x2_ASAP7_75t_R port map( A => n20, B => enable, Y => routing(6));
   U20 : NAND3xp33_ASAP7_75t_R port map( A => n1, B => n22, C => address(2), Y 
                           => n21);
   U21 : NAND3xp33_ASAP7_75t_R port map( A => n3, B => n4, C => enable, Y => 
                           n24);
   U3 : NOR2xp33_ASAP7_75t_R port map( A => n22, B => n23, Y => routing(4));
   U4 : NOR2xp33_ASAP7_75t_R port map( A => n23, B => n3, Y => routing(2));
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n21, B => n7, Y => routing(5));
   U6 : NOR2xp33_ASAP7_75t_R port map( A => address(0), B => address(1), Y => 
                           n20);
   U7 : NOR4xp25_ASAP7_75t_R port map( A => address(2), B => n20, C => n24, D 
                           => n2, Y => routing(3));
   U9 : NOR4xp25_ASAP7_75t_R port map( A => address(5), B => n23, C => n2, D =>
                           n4, Y => routing(1));
   U10 : NOR3xp33_ASAP7_75t_R port map( A => n5, B => address(1), C => n21, Y 
                           => routing(0));
   U12 : INVx1_ASAP7_75t_R port map( A => n24, Y => n1);
   U13 : INVx1_ASAP7_75t_R port map( A => address(4), Y => n2);
   U14 : INVx1_ASAP7_75t_R port map( A => address(5), Y => n3);
   U15 : INVx1_ASAP7_75t_R port map( A => address(3), Y => n4);
   U16 : INVx1_ASAP7_75t_R port map( A => address(0), Y => n5);
   U17 : INVx1_ASAP7_75t_R port map( A => n20, Y => n6);
   U18 : INVx1_ASAP7_75t_R port map( A => address(1), Y => n7);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT6_0 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (5 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (5 downto 0));

end rr_arbiter_no_delay_CNT6_0;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT6_0 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AO21x1_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI31xp33_ASAP7_75t_R
      port( A1, A2, A3, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OR3x1_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO32x1_ASAP7_75t_R
      port( A1, A2, A3, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_5_port, grant_4_port, grant_3_port, grant_2_port, grant_1_port,
      grant_0_port, pre_req_5_port, pre_req_4_port, pre_req_3_port, 
      pre_req_2_port, pre_req_1_port, pre_req_0_port, N2, N3, N4, N5, N6, 
      mask_pre_5_port, mask_pre_4_port, mask_pre_3_port, mask_pre_2_port, N20, 
      n6_port, n7, n14, n16, n18, n20_port, n22, n24, n1, n2_port, n3_port, 
      n4_port, n5_port, n8, n9, n10, n11, n12, n13, n15, n17, n19, n21, n23, 
      n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39
      , n40, n41, n42, n43, n44, n45, n46 : std_logic;

begin
   grant <= ( grant_5_port, grant_4_port, grant_3_port, grant_2_port, 
      grant_1_port, grant_0_port );
   
   U13 : AO32x1_ASAP7_75t_R port map( A1 => n6_port, A2 => req(5), A3 => 
                           n5_port, B1 => n15, B2 => mask_pre_5_port, Y => 
                           grant_5_port);
   U14 : AO32x1_ASAP7_75t_R port map( A1 => n6_port, A2 => req(4), A3 => n8, B1
                           => n17, B2 => mask_pre_4_port, Y => grant_4_port);
   U15 : AO32x1_ASAP7_75t_R port map( A1 => n6_port, A2 => req(3), A3 => n9, B1
                           => n19, B2 => mask_pre_3_port, Y => grant_3_port);
   U16 : AO32x1_ASAP7_75t_R port map( A1 => n6_port, A2 => req(2), A3 => n21, 
                           B1 => n10, B2 => mask_pre_2_port, Y => grant_2_port)
                           ;
   U20 : OR3x1_ASAP7_75t_R port map( A => mask_pre_3_port, B => mask_pre_5_port
                           , C => mask_pre_4_port, Y => n7);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_4_port, A2 => ack, B1 => 
                           grant_4_port, B2 => n46, Y => n14);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_3_port, A2 => ack, B1 => 
                           grant_3_port, B2 => n46, Y => n16);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_2_port, A2 => ack, B1 => 
                           grant_2_port, B2 => n46, Y => n18);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_5_port, A2 => ack, B1 => 
                           grant_5_port, B2 => n46, Y => n20_port);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n46, Y => n22);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n46, Y => n24);
   pre_req_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n18, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_2_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n22, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n24, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_0_port);
   pre_req_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n16, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_3_port);
   pre_req_reg_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n14, CLK => clk
                           , RESET => n25, SET => n23, QN => pre_req_4_port);
   pre_req_reg_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n20_port, CLK 
                           => clk, RESET => n25, SET => n23, QN => 
                           pre_req_5_port);
   U4 : TIELOx1_ASAP7_75t_R port map( L => n23);
   U5 : AND2x2_ASAP7_75t_R port map( A => n41, B => n39, Y => n1);
   U11 : AND2x2_ASAP7_75t_R port map( A => n42, B => n1, Y => n2_port);
   U12 : AND2x2_ASAP7_75t_R port map( A => n43, B => n2_port, Y => n3_port);
   U17 : AND2x2_ASAP7_75t_R port map( A => n44, B => n3_port, Y => n4_port);
   U18 : XOR2xp5_ASAP7_75t_R port map( A => n45, B => n4_port, Y => n5_port);
   U19 : XOR2xp5_ASAP7_75t_R port map( A => n44, B => n3_port, Y => n8);
   U21 : XOR2xp5_ASAP7_75t_R port map( A => n43, B => n2_port, Y => n9);
   U22 : XOR2xp5_ASAP7_75t_R port map( A => n36, B => n37, Y => n10);
   U23 : AND2x2_ASAP7_75t_R port map( A => n36, B => n37, Y => n11);
   U24 : AND2x2_ASAP7_75t_R port map( A => n35, B => n11, Y => n12);
   U25 : AND2x2_ASAP7_75t_R port map( A => n34, B => n12, Y => n13);
   U26 : XOR2xp5_ASAP7_75t_R port map( A => n33, B => n13, Y => n15);
   U27 : XOR2xp5_ASAP7_75t_R port map( A => n34, B => n12, Y => n17);
   U28 : XOR2xp5_ASAP7_75t_R port map( A => n35, B => n11, Y => n19);
   U29 : XOR2xp5_ASAP7_75t_R port map( A => n42, B => n1, Y => n21);
   U30 : NOR2xp33_ASAP7_75t_R port map( A => n40, B => n39, Y => grant_0_port);
   U31 : NOR3xp33_ASAP7_75t_R port map( A => n7, B => N20, C => mask_pre_2_port
                           , Y => n6_port);
   U32 : INVx1_ASAP7_75t_R port map( A => rst, Y => n25);
   U33 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_2_port, B => N3, C => n42,
                           Y => mask_pre_2_port);
   U34 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_1_port, B => N2, C => n41,
                           Y => N20);
   U35 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_3_port, B => N4, C => n43,
                           Y => mask_pre_3_port);
   U36 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_4_port, B => N5, C => n44,
                           Y => mask_pre_4_port);
   U37 : NOR3xp33_ASAP7_75t_R port map( A => pre_req_5_port, B => N6, C => n45,
                           Y => mask_pre_5_port);
   U38 : OAI31xp33_ASAP7_75t_R port map( A1 => n40, A2 => n38, A3 => n41, B => 
                           n37, Y => grant_1_port);
   U39 : XNOR2xp5_ASAP7_75t_R port map( A => n41, B => n39, Y => n38);
   U40 : NOR2xp33_ASAP7_75t_R port map( A => pre_req_1_port, B => 
                           pre_req_0_port, Y => n26);
   U41 : AO21x1_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => 
                           pre_req_1_port, B => n26, Y => N2);
   U42 : NOR2xp33_ASAP7_75t_R port map( A => n30, B => pre_req_2_port, Y => n27
                           );
   U43 : AO21x1_ASAP7_75t_R port map( A1 => n30, A2 => pre_req_2_port, B => n27
                           , Y => N3);
   U44 : NOR2xp33_ASAP7_75t_R port map( A => n31, B => pre_req_3_port, Y => n28
                           );
   U45 : AO21x1_ASAP7_75t_R port map( A1 => n31, A2 => pre_req_3_port, B => n28
                           , Y => N4);
   U46 : XNOR2xp5_ASAP7_75t_R port map( A => pre_req_4_port, B => n32, Y => N5)
                           ;
   U47 : NOR2xp33_ASAP7_75t_R port map( A => pre_req_4_port, B => n32, Y => n29
                           );
   U48 : XOR2xp5_ASAP7_75t_R port map( A => pre_req_5_port, B => n29, Y => N6);
   U49 : INVx1_ASAP7_75t_R port map( A => n26, Y => n30);
   U50 : INVx1_ASAP7_75t_R port map( A => n27, Y => n31);
   U51 : INVx1_ASAP7_75t_R port map( A => n28, Y => n32);
   U52 : INVx1_ASAP7_75t_R port map( A => mask_pre_5_port, Y => n33);
   U53 : INVx1_ASAP7_75t_R port map( A => mask_pre_4_port, Y => n34);
   U54 : INVx1_ASAP7_75t_R port map( A => mask_pre_3_port, Y => n35);
   U55 : INVx1_ASAP7_75t_R port map( A => mask_pre_2_port, Y => n36);
   U56 : INVx1_ASAP7_75t_R port map( A => N20, Y => n37);
   U57 : INVx1_ASAP7_75t_R port map( A => req(0), Y => n39);
   U58 : INVx1_ASAP7_75t_R port map( A => n6_port, Y => n40);
   U59 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n41);
   U60 : INVx1_ASAP7_75t_R port map( A => req(2), Y => n42);
   U61 : INVx1_ASAP7_75t_R port map( A => req(3), Y => n43);
   U62 : INVx1_ASAP7_75t_R port map( A => req(4), Y => n44);
   U63 : INVx1_ASAP7_75t_R port map( A => req(5), Y => n45);
   U64 : INVx1_ASAP7_75t_R port map( A => ack, Y => n46);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity seq_packet_counter_1_0 is

   port( clk, rst, allocated : in std_logic;  packet_len : in std_logic_vector 
         (3 downto 0);  enr_vc : in std_logic;  flit_count : out 
         std_logic_vector (3 downto 0));

end seq_packet_counter_1_0;

architecture SYN_rtl of seq_packet_counter_1_0 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI311xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, C1 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12 : std_logic;

begin
   flit_count <= ( flit_count_3_port, flit_count_2_port, flit_count_1_port, 
      flit_count_0_port );
   
   U11 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(3), B => n19, Y => n18)
                           ;
   U12 : NAND2xp5_ASAP7_75t_R port map( A => packet_len(2), B => n19, Y => n21)
                           ;
   U13 : OAI21xp5_ASAP7_75t_R port map( A1 => n19, A2 => n10, B => n22, Y => 
                           n20);
   U14 : NAND2xp5_ASAP7_75t_R port map( A => n23, B => n10, Y => n16);
   U15 : AOI21xp5_ASAP7_75t_R port map( A1 => n8, A2 => flit_count_0_port, B =>
                           n24, Y => n22);
   U26 : OAI311xp33_ASAP7_75t_R port map( A1 => n16, A2 => flit_count_3_port, 
                           A3 => flit_count_2_port, B1 => n17, C1 => n18, Y => 
                           n25);
   U27 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n8, B
                           => n20, C => flit_count_3_port, Y => n17);
   U28 : OAI221xp5_ASAP7_75t_R port map( A1 => flit_count_2_port, A2 => n16, B1
                           => n7, B2 => n11, C => n21, Y => n26);
   U29 : OAI221xp5_ASAP7_75t_R port map( A1 => n12, A2 => n8, B1 => n10, B2 => 
                           n22, C => n16, Y => n27);
   flit_count_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_0_port);
   flit_count_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_1_port);
   flit_count_int_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_2_port);
   flit_count_int_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n5, CLK 
                           => clk, RESET => n3, SET => n2, QN => 
                           flit_count_3_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n2);
   U4 : AOI221xp5_ASAP7_75t_R port map( A1 => packet_len(0), A2 => n19, B1 => 
                           n24, B2 => flit_count_0_port, C => n23, Y => n1);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n9, B => enr_vc, Y => n19);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => enr_vc, B => allocated, Y => n24);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n3);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => n19, B => flit_count_0_port, C => 
                           n24, Y => n23);
   U9 : INVx1_ASAP7_75t_R port map( A => n27, Y => n4);
   U10 : INVx1_ASAP7_75t_R port map( A => n25, Y => n5);
   U16 : INVx1_ASAP7_75t_R port map( A => n26, Y => n6);
   U17 : INVx1_ASAP7_75t_R port map( A => n20, Y => n7);
   U18 : INVx1_ASAP7_75t_R port map( A => n19, Y => n8);
   U19 : INVx1_ASAP7_75t_R port map( A => allocated, Y => n9);
   U20 : INVx1_ASAP7_75t_R port map( A => flit_count_1_port, Y => n10);
   U21 : INVx1_ASAP7_75t_R port map( A => flit_count_2_port, Y => n11);
   U22 : INVx1_ASAP7_75t_R port map( A => packet_len(1), Y => n12);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_0 is

   port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;  
         routing : out std_logic_vector (6 downto 0));

end routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_0;

architecture SYN_rtl of routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_0 is

   component dxyu_routing_Xis1_Yis1_Zis1_0
      port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;
            routing : out std_logic_vector (6 downto 0));
   end component;

begin
   
   dxyu_routing_1 : dxyu_routing_Xis1_Yis1_Zis1_0 port map( address(5) => 
                           address(5), address(4) => address(4), address(3) => 
                           address(3), address(2) => address(2), address(1) => 
                           address(1), address(0) => address(0), enable => 
                           enable, routing(6) => routing(6), routing(5) => 
                           routing(5), routing(4) => routing(4), routing(3) => 
                           routing(3), routing(2) => routing(2), routing(1) => 
                           routing(1), routing(0) => routing(0));

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity credit_count_single_vc_depth_out2_0 is

   port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
         std_logic);

end credit_count_single_vc_depth_out2_0;

architecture SYN_rtl of credit_count_single_vc_depth_out2_0 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_val_1_port, count_val_0_port, n12, n13, n14, n15, n16, n17, n1,
      n2, n3, n4, n5, n6 : std_logic;

begin
   
   U10 : NAND2xp5_ASAP7_75t_R port map( A => vc_write_tx, B => n17, Y => n16);
   U11 : NAND2xp5_ASAP7_75t_R port map( A => incr_rx, B => count_val_0_port, Y 
                           => n14);
   U15 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n5, A2 => n14, B => n15, C => 
                           n6, Y => n13);
   U16 : XNOR2xp5_ASAP7_75t_R port map( A => n14, B => n5, Y => n12);
   U17 : NAND3xp33_ASAP7_75t_R port map( A => n14, B => n6, C => n17, Y => 
                           credit_avail);
   U18 : XNOR2xp5_ASAP7_75t_R port map( A => count_val_0_port, B => incr_rx, Y 
                           => n17);
   count_val_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1, CLK => 
                           clk, RESET => n3, SET => n4, QN => count_val_1_port)
                           ;
   count_val_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2, CLK => 
                           clk, RESET => n4, SET => n3, QN => count_val_0_port)
                           ;
   U3 : TIELOx1_ASAP7_75t_R port map( L => n3);
   U4 : OA21x2_ASAP7_75t_R port map( A1 => n6, A2 => n12, B => n13, Y => n1);
   U5 : OA21x2_ASAP7_75t_R port map( A1 => vc_write_tx, A2 => n17, B => n16, Y 
                           => n2);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx, B => n14, Y => n15);
   U7 : INVx1_ASAP7_75t_R port map( A => rst, Y => n4);
   U8 : INVx1_ASAP7_75t_R port map( A => n16, Y => n5);
   U9 : INVx1_ASAP7_75t_R port map( A => count_val_1_port, Y => n6);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity rr_arbiter_no_delay_CNT2_0 is

   port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  ack
         : in std_logic;  grant : out std_logic_vector (1 downto 0));

end rr_arbiter_no_delay_CNT2_0;

architecture SYN_rr_arbiter_no_delay of rr_arbiter_no_delay_CNT2_0 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal grant_1_port, grant_0_port, pre_req_1_port, pre_req_0_port, n7, n9, 
      n11, n1, n2, n3, n4, n5 : std_logic;

begin
   grant <= ( grant_1_port, grant_0_port );
   
   U9 : AND2x2_ASAP7_75t_R port map( A => req(0), B => n7, Y => grant_0_port);
   U10 : NAND3xp33_ASAP7_75t_R port map( A => req(1), B => n5, C => 
                           pre_req_0_port, Y => n7);
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_1_port, A2 => ack, B1 => 
                           grant_1_port, B2 => n3, Y => n9);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => pre_req_0_port, A2 => ack, B1 => 
                           grant_0_port, B2 => n3, Y => n11);
   U7 : OAI21xp5_ASAP7_75t_R port map( A1 => req(0), A2 => n4, B => n7, Y => 
                           grant_1_port);
   pre_req_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n9, CLK => clk,
                           RESET => n2, SET => n1, QN => pre_req_1_port);
   pre_req_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n11, CLK => clk
                           , RESET => n2, SET => n1, QN => pre_req_0_port);
   U5 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U6 : INVx1_ASAP7_75t_R port map( A => rst, Y => n2);
   U8 : INVx1_ASAP7_75t_R port map( A => ack, Y => n3);
   U11 : INVx1_ASAP7_75t_R port map( A => req(1), Y => n4);
   U12 : INVx1_ASAP7_75t_R port map( A => pre_req_1_port, Y => n5);

end SYN_rr_arbiter_no_delay;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity header_arbiter_and_decoder_1_1_1_7_6_2_1_DXYU is

   port( clk, rst : in std_logic;  header : in std_logic_vector (19 downto 0); 
         valid_data_vc, enr_vc : in std_logic_vector (1 downto 0);  ack_vc : in
         std_logic;  granted_rq : out std_logic_vector (6 downto 0);  
         input_vc_in_use, packet_end, granted_vc : out std_logic_vector (1 
         downto 0));

end header_arbiter_and_decoder_1_1_1_7_6_2_1_DXYU;

architecture SYN_rtl of header_arbiter_and_decoder_1_1_1_7_6_2_1_DXYU is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVxp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component seq_packet_counter_1_1
      port( clk, rst, allocated : in std_logic;  packet_len : in 
            std_logic_vector (3 downto 0);  enr_vc : in std_logic;  flit_count 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component seq_packet_counter_1_2
      port( clk, rst, allocated : in std_logic;  packet_len : in 
            std_logic_vector (3 downto 0);  enr_vc : in std_logic;  flit_count 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_1
      port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;
            routing : out std_logic_vector (6 downto 0));
   end component;
   
   component rr_arbiter_no_delay_CNT2_1
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR5xp2_ASAP7_75t_R
      port( A, B, C, D, E : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic0_port, granted_rq_5_port, granted_rq_0, n14, 
      granted_vc_0_port, flit_count_values_1_3_port, flit_count_values_1_2_port
      , flit_count_values_1_1_port, flit_count_values_1_0_port, 
      flit_count_values_0_3_port, flit_count_values_0_2_port, 
      flit_count_values_0_1_port, flit_count_values_0_0_port, 
      new_package_vc_1_port, new_package_vc_0_port, 
      header_nxt_PACKET_LENGTH_3_port, header_nxt_PACKET_LENGTH_2_port, 
      header_nxt_PACKET_LENGTH_1_port, header_nxt_PACKET_LENGTH_0_port, 
      header_nxt_X_DEST_1_port, header_nxt_X_DEST_0_port, 
      header_nxt_Y_DEST_1_port, header_nxt_Y_DEST_0_port, 
      header_nxt_Z_DEST_1_port, header_nxt_Z_DEST_0_port, routing_en, 
      allocated_1_port, allocated_0_port, n10, n11, granted_vc_1_port, n2, n3, 
      n4, n5, n6, n8, n9, n12, n_1488, n_1489, n_1490, n_1491, n_1492 : 
      std_logic;

begin
   granted_rq <= ( X_Logic0_port, granted_rq_5_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, granted_rq_0 );
   granted_vc <= ( granted_vc_1_port, granted_vc_0_port );
   
   U2 : NAND2xp5_ASAP7_75t_R port map( A => n8, B => n9, Y => routing_en);
   U16 : NOR5xp2_ASAP7_75t_R port map( A => flit_count_values_1_2_port, B => 
                           flit_count_values_1_3_port, C => 
                           flit_count_values_1_1_port, D => n12, E => n3, Y => 
                           packet_end(1));
   U17 : NOR5xp2_ASAP7_75t_R port map( A => flit_count_values_0_2_port, B => 
                           flit_count_values_0_3_port, C => 
                           flit_count_values_0_1_port, D => n6, E => n5, Y => 
                           packet_end(0));
   U18 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc(1), B => n10, Y => 
                           new_package_vc_1_port);
   U19 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc(0), B => n11, Y => 
                           new_package_vc_0_port);
   U20 : AO22x1_ASAP7_75t_R port map( A1 => header(11), A2 => granted_vc_1_port
                           , B1 => header(1), B2 => n8, Y => 
                           header_nxt_Z_DEST_1_port);
   U21 : AO22x1_ASAP7_75t_R port map( A1 => header(10), A2 => granted_vc_1_port
                           , B1 => header(0), B2 => n8, Y => 
                           header_nxt_Z_DEST_0_port);
   U22 : AO22x1_ASAP7_75t_R port map( A1 => header(13), A2 => granted_vc_1_port
                           , B1 => header(3), B2 => n8, Y => 
                           header_nxt_Y_DEST_1_port);
   U23 : AO22x1_ASAP7_75t_R port map( A1 => header(12), A2 => granted_vc_1_port
                           , B1 => header(2), B2 => n8, Y => 
                           header_nxt_Y_DEST_0_port);
   U24 : AO22x1_ASAP7_75t_R port map( A1 => header(15), A2 => granted_vc_1_port
                           , B1 => header(5), B2 => n8, Y => 
                           header_nxt_X_DEST_1_port);
   U25 : AO22x1_ASAP7_75t_R port map( A1 => header(14), A2 => granted_vc_1_port
                           , B1 => header(4), B2 => n8, Y => 
                           header_nxt_X_DEST_0_port);
   U26 : AO22x1_ASAP7_75t_R port map( A1 => header(19), A2 => granted_vc_1_port
                           , B1 => header(9), B2 => n8, Y => 
                           header_nxt_PACKET_LENGTH_3_port);
   U27 : AO22x1_ASAP7_75t_R port map( A1 => header(18), A2 => granted_vc_1_port
                           , B1 => header(8), B2 => n8, Y => 
                           header_nxt_PACKET_LENGTH_2_port);
   U28 : AO22x1_ASAP7_75t_R port map( A1 => header(17), A2 => granted_vc_1_port
                           , B1 => header(7), B2 => n8, Y => 
                           header_nxt_PACKET_LENGTH_1_port);
   U29 : AO22x1_ASAP7_75t_R port map( A1 => header(16), A2 => granted_vc_1_port
                           , B1 => header(6), B2 => n8, Y => 
                           header_nxt_PACKET_LENGTH_0_port);
   rr_arbiter_no_delay_1 : rr_arbiter_no_delay_CNT2_1 port map( clk => clk, rst
                           => rst, req(1) => new_package_vc_1_port, req(0) => 
                           new_package_vc_0_port, ack => ack_vc, grant(1) => 
                           n14, grant(0) => granted_vc_0_port);
   routing_calc_1 : routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_1 port map( 
                           address(5) => header_nxt_X_DEST_1_port, address(4) 
                           => header_nxt_X_DEST_0_port, address(3) => 
                           header_nxt_Y_DEST_1_port, address(2) => 
                           header_nxt_Y_DEST_0_port, address(1) => 
                           header_nxt_Z_DEST_1_port, address(0) => 
                           header_nxt_Z_DEST_0_port, enable => routing_en, 
                           routing(6) => n_1488, routing(5) => 
                           granted_rq_5_port, routing(4) => n_1489, routing(3) 
                           => n_1490, routing(2) => n_1491, routing(1) => 
                           n_1492, routing(0) => granted_rq_0);
   seq_packet_counter_i_0 : seq_packet_counter_1_2 port map( clk => clk, rst =>
                           rst, allocated => allocated_0_port, packet_len(3) =>
                           header_nxt_PACKET_LENGTH_3_port, packet_len(2) => 
                           header_nxt_PACKET_LENGTH_2_port, packet_len(1) => 
                           header_nxt_PACKET_LENGTH_1_port, packet_len(0) => 
                           header_nxt_PACKET_LENGTH_0_port, enr_vc => enr_vc(0)
                           , flit_count(3) => flit_count_values_0_3_port, 
                           flit_count(2) => flit_count_values_0_2_port, 
                           flit_count(1) => flit_count_values_0_1_port, 
                           flit_count(0) => flit_count_values_0_0_port);
   seq_packet_counter_i_1 : seq_packet_counter_1_1 port map( clk => clk, rst =>
                           rst, allocated => allocated_1_port, packet_len(3) =>
                           header_nxt_PACKET_LENGTH_3_port, packet_len(2) => 
                           header_nxt_PACKET_LENGTH_2_port, packet_len(1) => 
                           header_nxt_PACKET_LENGTH_1_port, packet_len(0) => 
                           header_nxt_PACKET_LENGTH_0_port, enr_vc => n2, 
                           flit_count(3) => flit_count_values_1_3_port, 
                           flit_count(2) => flit_count_values_1_2_port, 
                           flit_count(1) => flit_count_values_1_1_port, 
                           flit_count(0) => flit_count_values_1_0_port);
   U3 : INVx1_ASAP7_75t_R port map( A => enr_vc(1), Y => n3);
   U4 : INVx1_ASAP7_75t_R port map( A => granted_vc_1_port, Y => n8);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n4, B => n9, Y => allocated_0_port)
                           ;
   U6 : NOR2xp33_ASAP7_75t_R port map( A => n8, B => n4, Y => allocated_1_port)
                           ;
   U7 : HB1xp67_ASAP7_75t_R port map( A => n14, Y => granted_vc_1_port);
   U8 : NOR4xp25_ASAP7_75t_R port map( A => flit_count_values_1_0_port, B => 
                           flit_count_values_1_1_port, C => 
                           flit_count_values_1_2_port, D => 
                           flit_count_values_1_3_port, Y => n10);
   U9 : NOR4xp25_ASAP7_75t_R port map( A => flit_count_values_0_0_port, B => 
                           flit_count_values_0_1_port, C => 
                           flit_count_values_0_2_port, D => 
                           flit_count_values_0_3_port, Y => n11);
   U10 : TIELOx1_ASAP7_75t_R port map( L => X_Logic0_port);
   U11 : INVxp67_ASAP7_75t_R port map( A => n3, Y => n2);
   U12 : INVx1_ASAP7_75t_R port map( A => ack_vc, Y => n4);
   U13 : INVx1_ASAP7_75t_R port map( A => enr_vc(0), Y => n5);
   U14 : INVx1_ASAP7_75t_R port map( A => flit_count_values_0_0_port, Y => n6);
   U15 : INVx1_ASAP7_75t_R port map( A => n11, Y => input_vc_in_use(0));
   U30 : INVx1_ASAP7_75t_R port map( A => granted_vc_0_port, Y => n9);
   U31 : INVx1_ASAP7_75t_R port map( A => flit_count_values_1_0_port, Y => n12)
                           ;
   U32 : INVx1_ASAP7_75t_R port map( A => n10, Y => input_vc_in_use(1));

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity header_arbiter_and_decoder_1_1_1_7_5_2_1_DXYU is

   port( clk, rst : in std_logic;  header : in std_logic_vector (19 downto 0); 
         valid_data_vc, enr_vc : in std_logic_vector (1 downto 0);  ack_vc : in
         std_logic;  granted_rq : out std_logic_vector (6 downto 0);  
         input_vc_in_use, packet_end, granted_vc : out std_logic_vector (1 
         downto 0));

end header_arbiter_and_decoder_1_1_1_7_5_2_1_DXYU;

architecture SYN_rtl of header_arbiter_and_decoder_1_1_1_7_5_2_1_DXYU is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component seq_packet_counter_1_3
      port( clk, rst, allocated : in std_logic;  packet_len : in 
            std_logic_vector (3 downto 0);  enr_vc : in std_logic;  flit_count 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component seq_packet_counter_1_4
      port( clk, rst, allocated : in std_logic;  packet_len : in 
            std_logic_vector (3 downto 0);  enr_vc : in std_logic;  flit_count 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_2
      port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;
            routing : out std_logic_vector (6 downto 0));
   end component;
   
   component rr_arbiter_no_delay_CNT2_2
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR5xp2_ASAP7_75t_R
      port( A, B, C, D, E : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n13, granted_vc_0_port, flit_count_values_1_3_port, 
      flit_count_values_1_2_port, flit_count_values_1_1_port, 
      flit_count_values_1_0_port, flit_count_values_0_3_port, 
      flit_count_values_0_2_port, flit_count_values_0_1_port, 
      flit_count_values_0_0_port, new_package_vc_1_port, new_package_vc_0_port,
      header_nxt_PACKET_LENGTH_3_port, header_nxt_PACKET_LENGTH_2_port, 
      header_nxt_PACKET_LENGTH_1_port, header_nxt_PACKET_LENGTH_0_port, 
      header_nxt_X_DEST_1_port, header_nxt_X_DEST_0_port, 
      header_nxt_Y_DEST_1_port, header_nxt_Y_DEST_0_port, 
      header_nxt_Z_DEST_1_port, header_nxt_Z_DEST_0_port, routing_en, 
      allocated_1_port, allocated_0_port, n10, n11, granted_vc_1_port, n2, n3, 
      n4, n5, n7, n8, n9, n_1493 : std_logic;

begin
   granted_vc <= ( granted_vc_1_port, granted_vc_0_port );
   
   U2 : NAND2xp5_ASAP7_75t_R port map( A => n7, B => n8, Y => routing_en);
   U16 : NOR5xp2_ASAP7_75t_R port map( A => flit_count_values_1_2_port, B => 
                           flit_count_values_1_3_port, C => 
                           flit_count_values_1_1_port, D => n9, E => n2, Y => 
                           packet_end(1));
   U17 : NOR5xp2_ASAP7_75t_R port map( A => flit_count_values_0_2_port, B => 
                           flit_count_values_0_3_port, C => 
                           flit_count_values_0_1_port, D => n5, E => n4, Y => 
                           packet_end(0));
   U18 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc(1), B => n10, Y => 
                           new_package_vc_1_port);
   U19 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc(0), B => n11, Y => 
                           new_package_vc_0_port);
   U20 : AO22x1_ASAP7_75t_R port map( A1 => header(11), A2 => granted_vc_1_port
                           , B1 => header(1), B2 => n7, Y => 
                           header_nxt_Z_DEST_1_port);
   U21 : AO22x1_ASAP7_75t_R port map( A1 => header(10), A2 => granted_vc_1_port
                           , B1 => header(0), B2 => n7, Y => 
                           header_nxt_Z_DEST_0_port);
   U22 : AO22x1_ASAP7_75t_R port map( A1 => header(13), A2 => granted_vc_1_port
                           , B1 => header(3), B2 => n7, Y => 
                           header_nxt_Y_DEST_1_port);
   U23 : AO22x1_ASAP7_75t_R port map( A1 => header(12), A2 => granted_vc_1_port
                           , B1 => header(2), B2 => n7, Y => 
                           header_nxt_Y_DEST_0_port);
   U24 : AO22x1_ASAP7_75t_R port map( A1 => header(15), A2 => granted_vc_1_port
                           , B1 => header(5), B2 => n7, Y => 
                           header_nxt_X_DEST_1_port);
   U25 : AO22x1_ASAP7_75t_R port map( A1 => header(14), A2 => granted_vc_1_port
                           , B1 => header(4), B2 => n7, Y => 
                           header_nxt_X_DEST_0_port);
   U26 : AO22x1_ASAP7_75t_R port map( A1 => header(19), A2 => granted_vc_1_port
                           , B1 => header(9), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_3_port);
   U27 : AO22x1_ASAP7_75t_R port map( A1 => header(18), A2 => granted_vc_1_port
                           , B1 => header(8), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_2_port);
   U28 : AO22x1_ASAP7_75t_R port map( A1 => header(17), A2 => granted_vc_1_port
                           , B1 => header(7), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_1_port);
   U29 : AO22x1_ASAP7_75t_R port map( A1 => header(16), A2 => granted_vc_1_port
                           , B1 => header(6), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_0_port);
   rr_arbiter_no_delay_1 : rr_arbiter_no_delay_CNT2_2 port map( clk => clk, rst
                           => rst, req(1) => new_package_vc_1_port, req(0) => 
                           new_package_vc_0_port, ack => ack_vc, grant(1) => 
                           n13, grant(0) => granted_vc_0_port);
   routing_calc_1 : routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_2 port map( 
                           address(5) => header_nxt_X_DEST_1_port, address(4) 
                           => header_nxt_X_DEST_0_port, address(3) => 
                           header_nxt_Y_DEST_1_port, address(2) => 
                           header_nxt_Y_DEST_0_port, address(1) => 
                           header_nxt_Z_DEST_1_port, address(0) => 
                           header_nxt_Z_DEST_0_port, enable => routing_en, 
                           routing(6) => granted_rq(6), routing(5) => n_1493, 
                           routing(4) => granted_rq(4), routing(3) => 
                           granted_rq(3), routing(2) => granted_rq(2), 
                           routing(1) => granted_rq(1), routing(0) => 
                           granted_rq(0));
   seq_packet_counter_i_0 : seq_packet_counter_1_4 port map( clk => clk, rst =>
                           rst, allocated => allocated_0_port, packet_len(3) =>
                           header_nxt_PACKET_LENGTH_3_port, packet_len(2) => 
                           header_nxt_PACKET_LENGTH_2_port, packet_len(1) => 
                           header_nxt_PACKET_LENGTH_1_port, packet_len(0) => 
                           header_nxt_PACKET_LENGTH_0_port, enr_vc => enr_vc(0)
                           , flit_count(3) => flit_count_values_0_3_port, 
                           flit_count(2) => flit_count_values_0_2_port, 
                           flit_count(1) => flit_count_values_0_1_port, 
                           flit_count(0) => flit_count_values_0_0_port);
   seq_packet_counter_i_1 : seq_packet_counter_1_3 port map( clk => clk, rst =>
                           rst, allocated => allocated_1_port, packet_len(3) =>
                           header_nxt_PACKET_LENGTH_3_port, packet_len(2) => 
                           header_nxt_PACKET_LENGTH_2_port, packet_len(1) => 
                           header_nxt_PACKET_LENGTH_1_port, packet_len(0) => 
                           header_nxt_PACKET_LENGTH_0_port, enr_vc => enr_vc(1)
                           , flit_count(3) => flit_count_values_1_3_port, 
                           flit_count(2) => flit_count_values_1_2_port, 
                           flit_count(1) => flit_count_values_1_1_port, 
                           flit_count(0) => flit_count_values_1_0_port);
   U3 : INVx1_ASAP7_75t_R port map( A => enr_vc(1), Y => n2);
   U4 : INVx1_ASAP7_75t_R port map( A => granted_vc_1_port, Y => n7);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n3, B => n8, Y => allocated_0_port)
                           ;
   U6 : NOR2xp33_ASAP7_75t_R port map( A => n7, B => n3, Y => allocated_1_port)
                           ;
   U7 : HB1xp67_ASAP7_75t_R port map( A => n13, Y => granted_vc_1_port);
   U8 : NOR4xp25_ASAP7_75t_R port map( A => flit_count_values_1_0_port, B => 
                           flit_count_values_1_1_port, C => 
                           flit_count_values_1_2_port, D => 
                           flit_count_values_1_3_port, Y => n10);
   U9 : NOR4xp25_ASAP7_75t_R port map( A => flit_count_values_0_0_port, B => 
                           flit_count_values_0_1_port, C => 
                           flit_count_values_0_2_port, D => 
                           flit_count_values_0_3_port, Y => n11);
   U10 : TIELOx1_ASAP7_75t_R port map( L => granted_rq(5));
   U11 : INVx1_ASAP7_75t_R port map( A => ack_vc, Y => n3);
   U12 : INVx1_ASAP7_75t_R port map( A => enr_vc(0), Y => n4);
   U13 : INVx1_ASAP7_75t_R port map( A => flit_count_values_0_0_port, Y => n5);
   U14 : INVx1_ASAP7_75t_R port map( A => n11, Y => input_vc_in_use(0));
   U15 : INVx1_ASAP7_75t_R port map( A => granted_vc_0_port, Y => n8);
   U30 : INVx1_ASAP7_75t_R port map( A => flit_count_values_1_0_port, Y => n9);
   U31 : INVx1_ASAP7_75t_R port map( A => n10, Y => input_vc_in_use(1));

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity header_arbiter_and_decoder_1_1_1_7_4_2_1_DXYU is

   port( clk, rst : in std_logic;  header : in std_logic_vector (19 downto 0); 
         valid_data_vc, enr_vc : in std_logic_vector (1 downto 0);  ack_vc : in
         std_logic;  granted_rq : out std_logic_vector (6 downto 0);  
         input_vc_in_use, packet_end, granted_vc : out std_logic_vector (1 
         downto 0));

end header_arbiter_and_decoder_1_1_1_7_4_2_1_DXYU;

architecture SYN_rtl of header_arbiter_and_decoder_1_1_1_7_4_2_1_DXYU is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component seq_packet_counter_1_5
      port( clk, rst, allocated : in std_logic;  packet_len : in 
            std_logic_vector (3 downto 0);  enr_vc : in std_logic;  flit_count 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component seq_packet_counter_1_6
      port( clk, rst, allocated : in std_logic;  packet_len : in 
            std_logic_vector (3 downto 0);  enr_vc : in std_logic;  flit_count 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_3
      port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;
            routing : out std_logic_vector (6 downto 0));
   end component;
   
   component rr_arbiter_no_delay_CNT2_3
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR5xp2_ASAP7_75t_R
      port( A, B, C, D, E : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic0_port, granted_rq_5, granted_rq_3_port, granted_rq_2_port, 
      granted_rq_1_port, granted_rq_0_port, n13, granted_vc_0_port, 
      flit_count_values_1_3_port, flit_count_values_1_2_port, 
      flit_count_values_1_1_port, flit_count_values_1_0_port, 
      flit_count_values_0_3_port, flit_count_values_0_2_port, 
      flit_count_values_0_1_port, flit_count_values_0_0_port, 
      new_package_vc_1_port, new_package_vc_0_port, 
      header_nxt_PACKET_LENGTH_3_port, header_nxt_PACKET_LENGTH_2_port, 
      header_nxt_PACKET_LENGTH_1_port, header_nxt_PACKET_LENGTH_0_port, 
      header_nxt_X_DEST_1_port, header_nxt_X_DEST_0_port, 
      header_nxt_Y_DEST_1_port, header_nxt_Y_DEST_0_port, 
      header_nxt_Z_DEST_1_port, header_nxt_Z_DEST_0_port, routing_en, 
      allocated_1_port, allocated_0_port, n10, n11, granted_vc_1_port, n2, n3, 
      n4, n5, n7, n8, n9, n_1494, n_1495 : std_logic;

begin
   granted_rq <= ( X_Logic0_port, granted_rq_5, X_Logic0_port, 
      granted_rq_3_port, granted_rq_2_port, granted_rq_1_port, 
      granted_rq_0_port );
   granted_vc <= ( granted_vc_1_port, granted_vc_0_port );
   
   U2 : NAND2xp5_ASAP7_75t_R port map( A => n7, B => n8, Y => routing_en);
   U16 : NOR5xp2_ASAP7_75t_R port map( A => flit_count_values_1_2_port, B => 
                           flit_count_values_1_3_port, C => 
                           flit_count_values_1_1_port, D => n9, E => n2, Y => 
                           packet_end(1));
   U17 : NOR5xp2_ASAP7_75t_R port map( A => flit_count_values_0_2_port, B => 
                           flit_count_values_0_3_port, C => 
                           flit_count_values_0_1_port, D => n5, E => n4, Y => 
                           packet_end(0));
   U18 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc(1), B => n10, Y => 
                           new_package_vc_1_port);
   U19 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc(0), B => n11, Y => 
                           new_package_vc_0_port);
   U20 : AO22x1_ASAP7_75t_R port map( A1 => header(11), A2 => granted_vc_1_port
                           , B1 => header(1), B2 => n7, Y => 
                           header_nxt_Z_DEST_1_port);
   U21 : AO22x1_ASAP7_75t_R port map( A1 => header(10), A2 => granted_vc_1_port
                           , B1 => header(0), B2 => n7, Y => 
                           header_nxt_Z_DEST_0_port);
   U22 : AO22x1_ASAP7_75t_R port map( A1 => header(13), A2 => granted_vc_1_port
                           , B1 => header(3), B2 => n7, Y => 
                           header_nxt_Y_DEST_1_port);
   U23 : AO22x1_ASAP7_75t_R port map( A1 => header(12), A2 => granted_vc_1_port
                           , B1 => header(2), B2 => n7, Y => 
                           header_nxt_Y_DEST_0_port);
   U24 : AO22x1_ASAP7_75t_R port map( A1 => header(15), A2 => granted_vc_1_port
                           , B1 => header(5), B2 => n7, Y => 
                           header_nxt_X_DEST_1_port);
   U25 : AO22x1_ASAP7_75t_R port map( A1 => header(14), A2 => granted_vc_1_port
                           , B1 => header(4), B2 => n7, Y => 
                           header_nxt_X_DEST_0_port);
   U26 : AO22x1_ASAP7_75t_R port map( A1 => header(19), A2 => granted_vc_1_port
                           , B1 => header(9), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_3_port);
   U27 : AO22x1_ASAP7_75t_R port map( A1 => header(18), A2 => granted_vc_1_port
                           , B1 => header(8), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_2_port);
   U28 : AO22x1_ASAP7_75t_R port map( A1 => header(17), A2 => granted_vc_1_port
                           , B1 => header(7), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_1_port);
   U29 : AO22x1_ASAP7_75t_R port map( A1 => header(16), A2 => granted_vc_1_port
                           , B1 => header(6), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_0_port);
   rr_arbiter_no_delay_1 : rr_arbiter_no_delay_CNT2_3 port map( clk => clk, rst
                           => rst, req(1) => new_package_vc_1_port, req(0) => 
                           new_package_vc_0_port, ack => ack_vc, grant(1) => 
                           n13, grant(0) => granted_vc_0_port);
   routing_calc_1 : routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_3 port map( 
                           address(5) => header_nxt_X_DEST_1_port, address(4) 
                           => header_nxt_X_DEST_0_port, address(3) => 
                           header_nxt_Y_DEST_1_port, address(2) => 
                           header_nxt_Y_DEST_0_port, address(1) => 
                           header_nxt_Z_DEST_1_port, address(0) => 
                           header_nxt_Z_DEST_0_port, enable => routing_en, 
                           routing(6) => n_1494, routing(5) => granted_rq_5, 
                           routing(4) => n_1495, routing(3) => 
                           granted_rq_3_port, routing(2) => granted_rq_2_port, 
                           routing(1) => granted_rq_1_port, routing(0) => 
                           granted_rq_0_port);
   seq_packet_counter_i_0 : seq_packet_counter_1_6 port map( clk => clk, rst =>
                           rst, allocated => allocated_0_port, packet_len(3) =>
                           header_nxt_PACKET_LENGTH_3_port, packet_len(2) => 
                           header_nxt_PACKET_LENGTH_2_port, packet_len(1) => 
                           header_nxt_PACKET_LENGTH_1_port, packet_len(0) => 
                           header_nxt_PACKET_LENGTH_0_port, enr_vc => enr_vc(0)
                           , flit_count(3) => flit_count_values_0_3_port, 
                           flit_count(2) => flit_count_values_0_2_port, 
                           flit_count(1) => flit_count_values_0_1_port, 
                           flit_count(0) => flit_count_values_0_0_port);
   seq_packet_counter_i_1 : seq_packet_counter_1_5 port map( clk => clk, rst =>
                           rst, allocated => allocated_1_port, packet_len(3) =>
                           header_nxt_PACKET_LENGTH_3_port, packet_len(2) => 
                           header_nxt_PACKET_LENGTH_2_port, packet_len(1) => 
                           header_nxt_PACKET_LENGTH_1_port, packet_len(0) => 
                           header_nxt_PACKET_LENGTH_0_port, enr_vc => enr_vc(1)
                           , flit_count(3) => flit_count_values_1_3_port, 
                           flit_count(2) => flit_count_values_1_2_port, 
                           flit_count(1) => flit_count_values_1_1_port, 
                           flit_count(0) => flit_count_values_1_0_port);
   U3 : INVx1_ASAP7_75t_R port map( A => enr_vc(1), Y => n2);
   U4 : NOR2xp33_ASAP7_75t_R port map( A => n3, B => n8, Y => allocated_0_port)
                           ;
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n7, B => n3, Y => allocated_1_port)
                           ;
   U6 : INVx1_ASAP7_75t_R port map( A => granted_vc_1_port, Y => n7);
   U7 : HB1xp67_ASAP7_75t_R port map( A => n13, Y => granted_vc_1_port);
   U8 : NOR4xp25_ASAP7_75t_R port map( A => flit_count_values_1_0_port, B => 
                           flit_count_values_1_1_port, C => 
                           flit_count_values_1_2_port, D => 
                           flit_count_values_1_3_port, Y => n10);
   U9 : NOR4xp25_ASAP7_75t_R port map( A => flit_count_values_0_0_port, B => 
                           flit_count_values_0_1_port, C => 
                           flit_count_values_0_2_port, D => 
                           flit_count_values_0_3_port, Y => n11);
   U10 : TIELOx1_ASAP7_75t_R port map( L => X_Logic0_port);
   U11 : INVx1_ASAP7_75t_R port map( A => ack_vc, Y => n3);
   U12 : INVx1_ASAP7_75t_R port map( A => enr_vc(0), Y => n4);
   U13 : INVx1_ASAP7_75t_R port map( A => flit_count_values_0_0_port, Y => n5);
   U14 : INVx1_ASAP7_75t_R port map( A => n11, Y => input_vc_in_use(0));
   U15 : INVx1_ASAP7_75t_R port map( A => granted_vc_0_port, Y => n8);
   U30 : INVx1_ASAP7_75t_R port map( A => flit_count_values_1_0_port, Y => n9);
   U31 : INVx1_ASAP7_75t_R port map( A => n10, Y => input_vc_in_use(1));

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity header_arbiter_and_decoder_1_1_1_7_3_2_1_DXYU is

   port( clk, rst : in std_logic;  header : in std_logic_vector (19 downto 0); 
         valid_data_vc, enr_vc : in std_logic_vector (1 downto 0);  ack_vc : in
         std_logic;  granted_rq : out std_logic_vector (6 downto 0);  
         input_vc_in_use, packet_end, granted_vc : out std_logic_vector (1 
         downto 0));

end header_arbiter_and_decoder_1_1_1_7_3_2_1_DXYU;

architecture SYN_rtl of header_arbiter_and_decoder_1_1_1_7_3_2_1_DXYU is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component seq_packet_counter_1_7
      port( clk, rst, allocated : in std_logic;  packet_len : in 
            std_logic_vector (3 downto 0);  enr_vc : in std_logic;  flit_count 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component seq_packet_counter_1_8
      port( clk, rst, allocated : in std_logic;  packet_len : in 
            std_logic_vector (3 downto 0);  enr_vc : in std_logic;  flit_count 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_4
      port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;
            routing : out std_logic_vector (6 downto 0));
   end component;
   
   component rr_arbiter_no_delay_CNT2_4
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR5xp2_ASAP7_75t_R
      port( A, B, C, D, E : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic0_port, granted_rq_5, granted_rq_1_port, granted_rq_0_port, 
      n13, granted_vc_0_port, flit_count_values_1_3_port, 
      flit_count_values_1_2_port, flit_count_values_1_1_port, 
      flit_count_values_1_0_port, flit_count_values_0_3_port, 
      flit_count_values_0_2_port, flit_count_values_0_1_port, 
      flit_count_values_0_0_port, new_package_vc_1_port, new_package_vc_0_port,
      header_nxt_PACKET_LENGTH_3_port, header_nxt_PACKET_LENGTH_2_port, 
      header_nxt_PACKET_LENGTH_1_port, header_nxt_PACKET_LENGTH_0_port, 
      header_nxt_X_DEST_1_port, header_nxt_X_DEST_0_port, 
      header_nxt_Y_DEST_1_port, header_nxt_Y_DEST_0_port, 
      header_nxt_Z_DEST_1_port, header_nxt_Z_DEST_0_port, routing_en, 
      allocated_1_port, allocated_0_port, n10, n11, granted_vc_1_port, n2, n3, 
      n4, n5, n7, n8, n9, n_1496, n_1497, n_1498, n_1499 : std_logic;

begin
   granted_rq <= ( X_Logic0_port, granted_rq_5, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, granted_rq_1_port, granted_rq_0_port );
   granted_vc <= ( granted_vc_1_port, granted_vc_0_port );
   
   U2 : NAND2xp5_ASAP7_75t_R port map( A => n7, B => n8, Y => routing_en);
   U16 : NOR5xp2_ASAP7_75t_R port map( A => flit_count_values_1_2_port, B => 
                           flit_count_values_1_3_port, C => 
                           flit_count_values_1_1_port, D => n9, E => n2, Y => 
                           packet_end(1));
   U17 : NOR5xp2_ASAP7_75t_R port map( A => flit_count_values_0_2_port, B => 
                           flit_count_values_0_3_port, C => 
                           flit_count_values_0_1_port, D => n5, E => n4, Y => 
                           packet_end(0));
   U18 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc(1), B => n10, Y => 
                           new_package_vc_1_port);
   U19 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc(0), B => n11, Y => 
                           new_package_vc_0_port);
   U20 : AO22x1_ASAP7_75t_R port map( A1 => header(11), A2 => granted_vc_1_port
                           , B1 => header(1), B2 => n7, Y => 
                           header_nxt_Z_DEST_1_port);
   U21 : AO22x1_ASAP7_75t_R port map( A1 => header(10), A2 => granted_vc_1_port
                           , B1 => header(0), B2 => n7, Y => 
                           header_nxt_Z_DEST_0_port);
   U22 : AO22x1_ASAP7_75t_R port map( A1 => header(13), A2 => granted_vc_1_port
                           , B1 => header(3), B2 => n7, Y => 
                           header_nxt_Y_DEST_1_port);
   U23 : AO22x1_ASAP7_75t_R port map( A1 => header(12), A2 => granted_vc_1_port
                           , B1 => header(2), B2 => n7, Y => 
                           header_nxt_Y_DEST_0_port);
   U24 : AO22x1_ASAP7_75t_R port map( A1 => header(15), A2 => granted_vc_1_port
                           , B1 => header(5), B2 => n7, Y => 
                           header_nxt_X_DEST_1_port);
   U25 : AO22x1_ASAP7_75t_R port map( A1 => header(14), A2 => granted_vc_1_port
                           , B1 => header(4), B2 => n7, Y => 
                           header_nxt_X_DEST_0_port);
   U26 : AO22x1_ASAP7_75t_R port map( A1 => header(19), A2 => granted_vc_1_port
                           , B1 => header(9), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_3_port);
   U27 : AO22x1_ASAP7_75t_R port map( A1 => header(18), A2 => granted_vc_1_port
                           , B1 => header(8), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_2_port);
   U28 : AO22x1_ASAP7_75t_R port map( A1 => header(17), A2 => granted_vc_1_port
                           , B1 => header(7), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_1_port);
   U29 : AO22x1_ASAP7_75t_R port map( A1 => header(16), A2 => granted_vc_1_port
                           , B1 => header(6), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_0_port);
   rr_arbiter_no_delay_1 : rr_arbiter_no_delay_CNT2_4 port map( clk => clk, rst
                           => rst, req(1) => new_package_vc_1_port, req(0) => 
                           new_package_vc_0_port, ack => ack_vc, grant(1) => 
                           n13, grant(0) => granted_vc_0_port);
   routing_calc_1 : routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_4 port map( 
                           address(5) => header_nxt_X_DEST_1_port, address(4) 
                           => header_nxt_X_DEST_0_port, address(3) => 
                           header_nxt_Y_DEST_1_port, address(2) => 
                           header_nxt_Y_DEST_0_port, address(1) => 
                           header_nxt_Z_DEST_1_port, address(0) => 
                           header_nxt_Z_DEST_0_port, enable => routing_en, 
                           routing(6) => n_1496, routing(5) => granted_rq_5, 
                           routing(4) => n_1497, routing(3) => n_1498, 
                           routing(2) => n_1499, routing(1) => 
                           granted_rq_1_port, routing(0) => granted_rq_0_port);
   seq_packet_counter_i_0 : seq_packet_counter_1_8 port map( clk => clk, rst =>
                           rst, allocated => allocated_0_port, packet_len(3) =>
                           header_nxt_PACKET_LENGTH_3_port, packet_len(2) => 
                           header_nxt_PACKET_LENGTH_2_port, packet_len(1) => 
                           header_nxt_PACKET_LENGTH_1_port, packet_len(0) => 
                           header_nxt_PACKET_LENGTH_0_port, enr_vc => enr_vc(0)
                           , flit_count(3) => flit_count_values_0_3_port, 
                           flit_count(2) => flit_count_values_0_2_port, 
                           flit_count(1) => flit_count_values_0_1_port, 
                           flit_count(0) => flit_count_values_0_0_port);
   seq_packet_counter_i_1 : seq_packet_counter_1_7 port map( clk => clk, rst =>
                           rst, allocated => allocated_1_port, packet_len(3) =>
                           header_nxt_PACKET_LENGTH_3_port, packet_len(2) => 
                           header_nxt_PACKET_LENGTH_2_port, packet_len(1) => 
                           header_nxt_PACKET_LENGTH_1_port, packet_len(0) => 
                           header_nxt_PACKET_LENGTH_0_port, enr_vc => enr_vc(1)
                           , flit_count(3) => flit_count_values_1_3_port, 
                           flit_count(2) => flit_count_values_1_2_port, 
                           flit_count(1) => flit_count_values_1_1_port, 
                           flit_count(0) => flit_count_values_1_0_port);
   U3 : INVx1_ASAP7_75t_R port map( A => enr_vc(1), Y => n2);
   U4 : INVx1_ASAP7_75t_R port map( A => granted_vc_1_port, Y => n7);
   U5 : HB1xp67_ASAP7_75t_R port map( A => n13, Y => granted_vc_1_port);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => n3, B => n8, Y => allocated_0_port)
                           ;
   U7 : NOR2xp33_ASAP7_75t_R port map( A => n7, B => n3, Y => allocated_1_port)
                           ;
   U8 : NOR4xp25_ASAP7_75t_R port map( A => flit_count_values_1_0_port, B => 
                           flit_count_values_1_1_port, C => 
                           flit_count_values_1_2_port, D => 
                           flit_count_values_1_3_port, Y => n10);
   U9 : NOR4xp25_ASAP7_75t_R port map( A => flit_count_values_0_0_port, B => 
                           flit_count_values_0_1_port, C => 
                           flit_count_values_0_2_port, D => 
                           flit_count_values_0_3_port, Y => n11);
   U10 : TIELOx1_ASAP7_75t_R port map( L => X_Logic0_port);
   U11 : INVx1_ASAP7_75t_R port map( A => ack_vc, Y => n3);
   U12 : INVx1_ASAP7_75t_R port map( A => enr_vc(0), Y => n4);
   U13 : INVx1_ASAP7_75t_R port map( A => flit_count_values_0_0_port, Y => n5);
   U14 : INVx1_ASAP7_75t_R port map( A => n11, Y => input_vc_in_use(0));
   U15 : INVx1_ASAP7_75t_R port map( A => granted_vc_0_port, Y => n8);
   U30 : INVx1_ASAP7_75t_R port map( A => flit_count_values_1_0_port, Y => n9);
   U31 : INVx1_ASAP7_75t_R port map( A => n10, Y => input_vc_in_use(1));

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity header_arbiter_and_decoder_1_1_1_7_2_2_1_DXYU is

   port( clk, rst : in std_logic;  header : in std_logic_vector (19 downto 0); 
         valid_data_vc, enr_vc : in std_logic_vector (1 downto 0);  ack_vc : in
         std_logic;  granted_rq : out std_logic_vector (6 downto 0);  
         input_vc_in_use, packet_end, granted_vc : out std_logic_vector (1 
         downto 0));

end header_arbiter_and_decoder_1_1_1_7_2_2_1_DXYU;

architecture SYN_rtl of header_arbiter_and_decoder_1_1_1_7_2_2_1_DXYU is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component seq_packet_counter_1_9
      port( clk, rst, allocated : in std_logic;  packet_len : in 
            std_logic_vector (3 downto 0);  enr_vc : in std_logic;  flit_count 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component seq_packet_counter_1_10
      port( clk, rst, allocated : in std_logic;  packet_len : in 
            std_logic_vector (3 downto 0);  enr_vc : in std_logic;  flit_count 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_5
      port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;
            routing : out std_logic_vector (6 downto 0));
   end component;
   
   component rr_arbiter_no_delay_CNT2_5
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR5xp2_ASAP7_75t_R
      port( A, B, C, D, E : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic0_port, granted_rq_5_port, granted_rq_4_port, 
      granted_rq_3_port, granted_rq_1, granted_rq_0, n13, granted_vc_0_port, 
      flit_count_values_1_3_port, flit_count_values_1_2_port, 
      flit_count_values_1_1_port, flit_count_values_1_0_port, 
      flit_count_values_0_3_port, flit_count_values_0_2_port, 
      flit_count_values_0_1_port, flit_count_values_0_0_port, 
      new_package_vc_1_port, new_package_vc_0_port, 
      header_nxt_PACKET_LENGTH_3_port, header_nxt_PACKET_LENGTH_2_port, 
      header_nxt_PACKET_LENGTH_1_port, header_nxt_PACKET_LENGTH_0_port, 
      header_nxt_X_DEST_1_port, header_nxt_X_DEST_0_port, 
      header_nxt_Y_DEST_1_port, header_nxt_Y_DEST_0_port, 
      header_nxt_Z_DEST_1_port, header_nxt_Z_DEST_0_port, routing_en, 
      allocated_1_port, allocated_0_port, n10, n11, granted_vc_1_port, n2, n3, 
      n4, n5, n7, n8, n9, n_1500, n_1501 : std_logic;

begin
   granted_rq <= ( X_Logic0_port, granted_rq_5_port, granted_rq_4_port, 
      granted_rq_3_port, X_Logic0_port, granted_rq_1, granted_rq_0 );
   granted_vc <= ( granted_vc_1_port, granted_vc_0_port );
   
   U2 : NAND2xp5_ASAP7_75t_R port map( A => n7, B => n8, Y => routing_en);
   U16 : NOR5xp2_ASAP7_75t_R port map( A => flit_count_values_1_2_port, B => 
                           flit_count_values_1_3_port, C => 
                           flit_count_values_1_1_port, D => n9, E => n2, Y => 
                           packet_end(1));
   U17 : NOR5xp2_ASAP7_75t_R port map( A => flit_count_values_0_2_port, B => 
                           flit_count_values_0_3_port, C => 
                           flit_count_values_0_1_port, D => n5, E => n4, Y => 
                           packet_end(0));
   U18 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc(1), B => n10, Y => 
                           new_package_vc_1_port);
   U19 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc(0), B => n11, Y => 
                           new_package_vc_0_port);
   U20 : AO22x1_ASAP7_75t_R port map( A1 => header(11), A2 => granted_vc_1_port
                           , B1 => header(1), B2 => n7, Y => 
                           header_nxt_Z_DEST_1_port);
   U21 : AO22x1_ASAP7_75t_R port map( A1 => header(10), A2 => granted_vc_1_port
                           , B1 => header(0), B2 => n7, Y => 
                           header_nxt_Z_DEST_0_port);
   U22 : AO22x1_ASAP7_75t_R port map( A1 => header(13), A2 => granted_vc_1_port
                           , B1 => header(3), B2 => n7, Y => 
                           header_nxt_Y_DEST_1_port);
   U23 : AO22x1_ASAP7_75t_R port map( A1 => header(12), A2 => granted_vc_1_port
                           , B1 => header(2), B2 => n7, Y => 
                           header_nxt_Y_DEST_0_port);
   U24 : AO22x1_ASAP7_75t_R port map( A1 => header(15), A2 => granted_vc_1_port
                           , B1 => header(5), B2 => n7, Y => 
                           header_nxt_X_DEST_1_port);
   U25 : AO22x1_ASAP7_75t_R port map( A1 => header(14), A2 => granted_vc_1_port
                           , B1 => header(4), B2 => n7, Y => 
                           header_nxt_X_DEST_0_port);
   U26 : AO22x1_ASAP7_75t_R port map( A1 => header(19), A2 => granted_vc_1_port
                           , B1 => header(9), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_3_port);
   U27 : AO22x1_ASAP7_75t_R port map( A1 => header(18), A2 => granted_vc_1_port
                           , B1 => header(8), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_2_port);
   U28 : AO22x1_ASAP7_75t_R port map( A1 => header(17), A2 => granted_vc_1_port
                           , B1 => header(7), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_1_port);
   U29 : AO22x1_ASAP7_75t_R port map( A1 => header(16), A2 => granted_vc_1_port
                           , B1 => header(6), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_0_port);
   rr_arbiter_no_delay_1 : rr_arbiter_no_delay_CNT2_5 port map( clk => clk, rst
                           => rst, req(1) => new_package_vc_1_port, req(0) => 
                           new_package_vc_0_port, ack => ack_vc, grant(1) => 
                           n13, grant(0) => granted_vc_0_port);
   routing_calc_1 : routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_5 port map( 
                           address(5) => header_nxt_X_DEST_1_port, address(4) 
                           => header_nxt_X_DEST_0_port, address(3) => 
                           header_nxt_Y_DEST_1_port, address(2) => 
                           header_nxt_Y_DEST_0_port, address(1) => 
                           header_nxt_Z_DEST_1_port, address(0) => 
                           header_nxt_Z_DEST_0_port, enable => routing_en, 
                           routing(6) => n_1500, routing(5) => 
                           granted_rq_5_port, routing(4) => granted_rq_4_port, 
                           routing(3) => granted_rq_3_port, routing(2) => 
                           n_1501, routing(1) => granted_rq_1, routing(0) => 
                           granted_rq_0);
   seq_packet_counter_i_0 : seq_packet_counter_1_10 port map( clk => clk, rst 
                           => rst, allocated => allocated_0_port, packet_len(3)
                           => header_nxt_PACKET_LENGTH_3_port, packet_len(2) =>
                           header_nxt_PACKET_LENGTH_2_port, packet_len(1) => 
                           header_nxt_PACKET_LENGTH_1_port, packet_len(0) => 
                           header_nxt_PACKET_LENGTH_0_port, enr_vc => enr_vc(0)
                           , flit_count(3) => flit_count_values_0_3_port, 
                           flit_count(2) => flit_count_values_0_2_port, 
                           flit_count(1) => flit_count_values_0_1_port, 
                           flit_count(0) => flit_count_values_0_0_port);
   seq_packet_counter_i_1 : seq_packet_counter_1_9 port map( clk => clk, rst =>
                           rst, allocated => allocated_1_port, packet_len(3) =>
                           header_nxt_PACKET_LENGTH_3_port, packet_len(2) => 
                           header_nxt_PACKET_LENGTH_2_port, packet_len(1) => 
                           header_nxt_PACKET_LENGTH_1_port, packet_len(0) => 
                           header_nxt_PACKET_LENGTH_0_port, enr_vc => enr_vc(1)
                           , flit_count(3) => flit_count_values_1_3_port, 
                           flit_count(2) => flit_count_values_1_2_port, 
                           flit_count(1) => flit_count_values_1_1_port, 
                           flit_count(0) => flit_count_values_1_0_port);
   U3 : INVx1_ASAP7_75t_R port map( A => enr_vc(1), Y => n2);
   U4 : INVx1_ASAP7_75t_R port map( A => granted_vc_1_port, Y => n7);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n3, B => n8, Y => allocated_0_port)
                           ;
   U6 : NOR2xp33_ASAP7_75t_R port map( A => n7, B => n3, Y => allocated_1_port)
                           ;
   U7 : HB1xp67_ASAP7_75t_R port map( A => n13, Y => granted_vc_1_port);
   U8 : NOR4xp25_ASAP7_75t_R port map( A => flit_count_values_1_0_port, B => 
                           flit_count_values_1_1_port, C => 
                           flit_count_values_1_2_port, D => 
                           flit_count_values_1_3_port, Y => n10);
   U9 : NOR4xp25_ASAP7_75t_R port map( A => flit_count_values_0_0_port, B => 
                           flit_count_values_0_1_port, C => 
                           flit_count_values_0_2_port, D => 
                           flit_count_values_0_3_port, Y => n11);
   U10 : TIELOx1_ASAP7_75t_R port map( L => X_Logic0_port);
   U11 : INVx1_ASAP7_75t_R port map( A => ack_vc, Y => n3);
   U12 : INVx1_ASAP7_75t_R port map( A => enr_vc(0), Y => n4);
   U13 : INVx1_ASAP7_75t_R port map( A => flit_count_values_0_0_port, Y => n5);
   U14 : INVx1_ASAP7_75t_R port map( A => n11, Y => input_vc_in_use(0));
   U15 : INVx1_ASAP7_75t_R port map( A => granted_vc_0_port, Y => n8);
   U30 : INVx1_ASAP7_75t_R port map( A => flit_count_values_1_0_port, Y => n9);
   U31 : INVx1_ASAP7_75t_R port map( A => n10, Y => input_vc_in_use(1));

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity vc_output_allocator_port_num7_vc_num_out2_0 is

   port( clk, rst : in std_logic;  rq_vc_out : in std_logic_vector (5 downto 0)
         ;  granted_vc, packet_end : in std_logic_vector (11 downto 0);  
         crossbar_ctrl_vec : out std_logic_vector (5 downto 0);  vc_sel_enc, 
         output_vc_in_use : out std_logic_vector (1 downto 0);  ack_rq_vc_out :
         out std_logic_vector (5 downto 0));

end vc_output_allocator_port_num7_vc_num_out2_0;

architecture SYN_rtl of vc_output_allocator_port_num7_vc_num_out2_0 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OA21x2_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21xp5_ASAP7_75t_R
      port( A1, A2, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component rr_arbiter_no_delay_CNT6_6
      port( clk, rst : in std_logic;  req : in std_logic_vector (5 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (5 downto 0));
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI211xp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OA211x2_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1O1Ixp25_ASAP7_75t_R
      port( A1, A2, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal crossbar_ctrl_vec_5_port, crossbar_ctrl_vec_4_port, n33, 
      crossbar_ctrl_vec_2_port, crossbar_ctrl_vec_1_port, n34, 
      vc_sel_enc_1_0_port, vc_sel_enc_0_0_port, output_vc_in_use_1_port, 
      output_vc_in_use_0_port, vc_available, grant_5_port, grant_4_port, 
      grant_3_port, grant_2_port, grant_1_port, grant_0_port, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n87
      , n88, n91, n1, n2, n3, n4, n5, crossbar_ctrl_vec_3_port, 
      crossbar_ctrl_vec_0_port, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      : std_logic;

begin
   crossbar_ctrl_vec <= ( crossbar_ctrl_vec_5_port, crossbar_ctrl_vec_4_port, 
      crossbar_ctrl_vec_3_port, crossbar_ctrl_vec_2_port, 
      crossbar_ctrl_vec_1_port, crossbar_ctrl_vec_0_port );
   vc_sel_enc <= ( vc_sel_enc_1_0_port, vc_sel_enc_0_0_port );
   output_vc_in_use <= ( output_vc_in_use_1_port, output_vc_in_use_0_port );
   
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => n40, A2 => n13, B1 => n41, B2 => 
                           n28, Y => n83);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => n42, A2 => n13, B1 => n41, B2 => 
                           n29, Y => n84);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => n43, A2 => n13, B1 => n41, B2 => 
                           n30, Y => n85);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => n40, A2 => n16, B1 => n44, B2 => 
                           n24, Y => n87);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => n42, A2 => n16, B1 => n44, B2 => 
                           n25, Y => n88);
   U28 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n47, A2 => n48, B => n26, C => 
                           n49, Y => n46);
   U30 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n23, B => n53, C => vc_sel_enc_0_0_port, Y => n52);
   U31 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(2), B => 
                           crossbar_ctrl_vec_0_port, Y => n53);
   U33 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n31, B => n54, C => n25, Y => n48);
   U34 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(10), B => 
                           crossbar_ctrl_vec_0_port, Y => n54);
   U35 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n21, B => n55, C => n24, Y => n47);
   U36 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(6), B => 
                           crossbar_ctrl_vec_0_port, Y => n55);
   U37 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n56, A2 => n57, B => 
                           vc_sel_enc_0_0_port, C => n27, Y => n45);
   U38 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n32, B => n58, C => n25, Y => n57);
   U39 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(11), B => 
                           crossbar_ctrl_vec_0_port, Y => n58);
   U40 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_0_port, A2 =>
                           n20, B => n59, C => n24, Y => n56);
   U41 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(7), B => 
                           crossbar_ctrl_vec_0_port, Y => n59);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => n43, A2 => n16, B1 => n44, B2 => 
                           n26, Y => n91);
   U52 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_3_port, A2 =>
                           n22, B => n79, C => n30, Y => n78);
   U53 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(3), B => 
                           crossbar_ctrl_vec_3_port, Y => n79);
   U54 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec_3_port, A2 =>
                           n23, B => n80, C => vc_sel_enc_1_0_port, Y => n77);
   U55 : NAND2xp5_ASAP7_75t_R port map( A => packet_end(2), B => 
                           crossbar_ctrl_vec_3_port, Y => n80);
   U58 : NAND2xp5_ASAP7_75t_R port map( A => output_vc_in_use_1_port, B => 
                           output_vc_in_use_0_port, Y => vc_available);
   U81 : A2O1A1O1Ixp25_ASAP7_75t_R port map( A1 => packet_end(3), A2 => 
                           crossbar_ctrl_vec_0_port, B => n51, C => 
                           vc_sel_enc_0_0_port, D => n52, Y => n50);
   U82 : OA211x2_ASAP7_75t_R port map( A1 => n19, A2 => n61, B => n62, C => n63
                           , Y => n43);
   U83 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(9), A2 => n64, B =>
                           n65, C => n18, Y => n63);
   U84 : AND2x2_ASAP7_75t_R port map( A => granted_vc(11), B => n17, Y => n65);
   U85 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(5), A2 => n64, B =>
                           n66, C => n19, Y => n62);
   U86 : AND2x2_ASAP7_75t_R port map( A => granted_vc(7), B => n17, Y => n66);
   U87 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(1), A2 => n64, B =>
                           n67, C => n42, Y => n61);
   U88 : AND2x2_ASAP7_75t_R port map( A => granted_vc(3), B => n17, Y => n67);
   U89 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n70, A2 => n71, B => n30, C =>
                           output_vc_in_use_1_port, Y => n69);
   U90 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(7), A2 => 
                           crossbar_ctrl_vec_3_port, B => n72, C => 
                           crossbar_ctrl_vec_4_port, Y => n71);
   U91 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(11), A2 => 
                           crossbar_ctrl_vec_3_port, B => n73, C => 
                           crossbar_ctrl_vec_5_port, Y => n70);
   U92 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n74, A2 => n75, B => 
                           vc_sel_enc_1_0_port, C => n76, Y => n68);
   U93 : OAI211xp5_ASAP7_75t_R port map( A1 => n77, A2 => n78, B => n28, C => 
                           n29, Y => n76);
   U94 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(6), A2 => 
                           crossbar_ctrl_vec_3_port, B => n81, C => 
                           crossbar_ctrl_vec_4_port, Y => n75);
   U95 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(10), A2 => 
                           crossbar_ctrl_vec_3_port, B => n82, C => 
                           crossbar_ctrl_vec_5_port, Y => n74);
   U96 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_5_port, Y 
                           => ack_rq_vc_out(5));
   U97 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_4_port, Y 
                           => ack_rq_vc_out(4));
   U98 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_3_port, Y 
                           => ack_rq_vc_out(3));
   U99 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_2_port, Y 
                           => ack_rq_vc_out(2));
   U100 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_1_port, Y 
                           => ack_rq_vc_out(1));
   U101 : AND2x2_ASAP7_75t_R port map( A => vc_available, B => grant_0_port, Y 
                           => ack_rq_vc_out(0));
   rr_arbiter : rr_arbiter_no_delay_CNT6_6 port map( clk => clk, rst => rst, 
                           req(5) => rq_vc_out(5), req(4) => rq_vc_out(4), 
                           req(3) => rq_vc_out(3), req(2) => rq_vc_out(2), 
                           req(1) => rq_vc_out(1), req(0) => rq_vc_out(0), ack 
                           => vc_available, grant(5) => grant_5_port, grant(4) 
                           => grant_4_port, grant(3) => grant_3_port, grant(2) 
                           => grant_2_port, grant(1) => grant_1_port, grant(0) 
                           => grant_0_port);
   vc_sel_enc_int_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n10, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           vc_sel_enc_1_0_port);
   crossbar_sels_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n11, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_4_port);
   crossbar_sels_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n12, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_5_port);
   crossbar_sels_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK
                           => clk, RESET => n8, SET => n5, QN => n33);
   vc_sel_enc_int_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n9, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           vc_sel_enc_0_0_port);
   crossbar_sels_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n15, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_2_port);
   crossbar_sels_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n14, 
                           CLK => clk, RESET => n8, SET => n5, QN => 
                           crossbar_ctrl_vec_1_port);
   crossbar_sels_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n3, CLK
                           => clk, RESET => n8, SET => n5, QN => n34);
   output_vc_in_use_int_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2
                           , CLK => clk, RESET => n8, SET => n5, QN => 
                           output_vc_in_use_1_port);
   output_vc_in_use_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n1
                           , CLK => clk, RESET => n8, SET => n5, QN => 
                           output_vc_in_use_0_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n5);
   U4 : AOI21xp5_ASAP7_75t_R port map( A1 => n45, A2 => n46, B => n44, Y => n1)
                           ;
   U5 : OA21x2_ASAP7_75t_R port map( A1 => n68, A2 => n69, B => n13, Y => n2);
   U6 : AOI22xp5_ASAP7_75t_R port map( A1 => n17, A2 => n44, B1 => n16, B2 => 
                           crossbar_ctrl_vec_0_port, Y => n3);
   U7 : AOI22xp5_ASAP7_75t_R port map( A1 => n17, A2 => n41, B1 => n13, B2 => 
                           crossbar_ctrl_vec_3_port, Y => n4);
   U8 : NOR3xp33_ASAP7_75t_R port map( A => grant_3_port, B => grant_5_port, C 
                           => grant_1_port, Y => n64);
   U9 : NOR2xp33_ASAP7_75t_R port map( A => grant_3_port, B => grant_2_port, Y 
                           => n40);
   U10 : NOR4xp25_ASAP7_75t_R port map( A => n17, B => grant_0_port, C => 
                           grant_2_port, D => grant_4_port, Y => n60);
   U11 : NOR2xp33_ASAP7_75t_R port map( A => grant_5_port, B => grant_4_port, Y
                           => n42);
   U12 : INVx1_ASAP7_75t_R port map( A => rst, Y => n8);
   U13 : NOR3xp33_ASAP7_75t_R port map( A => n50, B => crossbar_ctrl_vec_2_port
                           , C => crossbar_ctrl_vec_1_port, Y => n49);
   U14 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_0_port, B => n22
                           , Y => n51);
   U15 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n20
                           , Y => n72);
   U16 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n21
                           , Y => n81);
   U17 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n31
                           , Y => n82);
   U18 : HB1xp67_ASAP7_75t_R port map( A => n33, Y => crossbar_ctrl_vec_3_port)
                           ;
   U19 : HB1xp67_ASAP7_75t_R port map( A => n34, Y => crossbar_ctrl_vec_0_port)
                           ;
   U20 : NOR2xp33_ASAP7_75t_R port map( A => n60, B => output_vc_in_use_0_port,
                           Y => n44);
   U21 : NOR3xp33_ASAP7_75t_R port map( A => n60, B => output_vc_in_use_1_port,
                           C => n27, Y => n41);
   U22 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec_3_port, B => n32
                           , Y => n73);
   U29 : INVx1_ASAP7_75t_R port map( A => n91, Y => n9);
   U32 : INVx1_ASAP7_75t_R port map( A => n85, Y => n10);
   U43 : INVx1_ASAP7_75t_R port map( A => n83, Y => n11);
   U44 : INVx1_ASAP7_75t_R port map( A => n84, Y => n12);
   U45 : INVx1_ASAP7_75t_R port map( A => n41, Y => n13);
   U46 : INVx1_ASAP7_75t_R port map( A => n87, Y => n14);
   U47 : INVx1_ASAP7_75t_R port map( A => n88, Y => n15);
   U48 : INVx1_ASAP7_75t_R port map( A => n44, Y => n16);
   U49 : INVx1_ASAP7_75t_R port map( A => n64, Y => n17);
   U50 : INVx1_ASAP7_75t_R port map( A => n42, Y => n18);
   U51 : INVx1_ASAP7_75t_R port map( A => n40, Y => n19);
   U56 : INVx1_ASAP7_75t_R port map( A => packet_end(5), Y => n20);
   U57 : INVx1_ASAP7_75t_R port map( A => packet_end(4), Y => n21);
   U59 : INVx1_ASAP7_75t_R port map( A => packet_end(1), Y => n22);
   U60 : INVx1_ASAP7_75t_R port map( A => packet_end(0), Y => n23);
   U61 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_1_port, Y => n24);
   U62 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_2_port, Y => n25);
   U63 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_0_0_port, Y => n26);
   U64 : INVx1_ASAP7_75t_R port map( A => output_vc_in_use_0_port, Y => n27);
   U65 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_4_port, Y => n28);
   U66 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_5_port, Y => n29);
   U67 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_1_0_port, Y => n30);
   U68 : INVx1_ASAP7_75t_R port map( A => packet_end(8), Y => n31);
   U69 : INVx1_ASAP7_75t_R port map( A => packet_end(9), Y => n32);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity header_arbiter_and_decoder_1_1_1_7_1_2_1_DXYU is

   port( clk, rst : in std_logic;  header : in std_logic_vector (19 downto 0); 
         valid_data_vc, enr_vc : in std_logic_vector (1 downto 0);  ack_vc : in
         std_logic;  granted_rq : out std_logic_vector (6 downto 0);  
         input_vc_in_use, packet_end, granted_vc : out std_logic_vector (1 
         downto 0));

end header_arbiter_and_decoder_1_1_1_7_1_2_1_DXYU;

architecture SYN_rtl of header_arbiter_and_decoder_1_1_1_7_1_2_1_DXYU is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component seq_packet_counter_1_11
      port( clk, rst, allocated : in std_logic;  packet_len : in 
            std_logic_vector (3 downto 0);  enr_vc : in std_logic;  flit_count 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component seq_packet_counter_1_12
      port( clk, rst, allocated : in std_logic;  packet_len : in 
            std_logic_vector (3 downto 0);  enr_vc : in std_logic;  flit_count 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_6
      port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;
            routing : out std_logic_vector (6 downto 0));
   end component;
   
   component rr_arbiter_no_delay_CNT2_6
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR5xp2_ASAP7_75t_R
      port( A, B, C, D, E : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic0_port, granted_rq_5_port, granted_rq_3, granted_rq_0, n13, 
      granted_vc_0_port, flit_count_values_1_3_port, flit_count_values_1_2_port
      , flit_count_values_1_1_port, flit_count_values_1_0_port, 
      flit_count_values_0_3_port, flit_count_values_0_2_port, 
      flit_count_values_0_1_port, flit_count_values_0_0_port, 
      new_package_vc_1_port, new_package_vc_0_port, 
      header_nxt_PACKET_LENGTH_3_port, header_nxt_PACKET_LENGTH_2_port, 
      header_nxt_PACKET_LENGTH_1_port, header_nxt_PACKET_LENGTH_0_port, 
      header_nxt_X_DEST_1_port, header_nxt_X_DEST_0_port, 
      header_nxt_Y_DEST_1_port, header_nxt_Y_DEST_0_port, 
      header_nxt_Z_DEST_1_port, header_nxt_Z_DEST_0_port, routing_en, 
      allocated_1_port, allocated_0_port, n10, n11, granted_vc_1_port, n2, n3, 
      n4, n5, n7, n8, n9, n_1502, n_1503, n_1504, n_1505 : std_logic;

begin
   granted_rq <= ( X_Logic0_port, granted_rq_5_port, X_Logic0_port, 
      granted_rq_3, X_Logic0_port, X_Logic0_port, granted_rq_0 );
   granted_vc <= ( granted_vc_1_port, granted_vc_0_port );
   
   U2 : NAND2xp5_ASAP7_75t_R port map( A => n7, B => n8, Y => routing_en);
   U16 : NOR5xp2_ASAP7_75t_R port map( A => flit_count_values_1_2_port, B => 
                           flit_count_values_1_3_port, C => 
                           flit_count_values_1_1_port, D => n9, E => n2, Y => 
                           packet_end(1));
   U17 : NOR5xp2_ASAP7_75t_R port map( A => flit_count_values_0_2_port, B => 
                           flit_count_values_0_3_port, C => 
                           flit_count_values_0_1_port, D => n5, E => n4, Y => 
                           packet_end(0));
   U18 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc(1), B => n10, Y => 
                           new_package_vc_1_port);
   U19 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc(0), B => n11, Y => 
                           new_package_vc_0_port);
   U20 : AO22x1_ASAP7_75t_R port map( A1 => header(11), A2 => granted_vc_1_port
                           , B1 => header(1), B2 => n7, Y => 
                           header_nxt_Z_DEST_1_port);
   U21 : AO22x1_ASAP7_75t_R port map( A1 => header(10), A2 => granted_vc_1_port
                           , B1 => header(0), B2 => n7, Y => 
                           header_nxt_Z_DEST_0_port);
   U22 : AO22x1_ASAP7_75t_R port map( A1 => header(13), A2 => granted_vc_1_port
                           , B1 => header(3), B2 => n7, Y => 
                           header_nxt_Y_DEST_1_port);
   U23 : AO22x1_ASAP7_75t_R port map( A1 => header(12), A2 => granted_vc_1_port
                           , B1 => header(2), B2 => n7, Y => 
                           header_nxt_Y_DEST_0_port);
   U24 : AO22x1_ASAP7_75t_R port map( A1 => header(15), A2 => granted_vc_1_port
                           , B1 => header(5), B2 => n7, Y => 
                           header_nxt_X_DEST_1_port);
   U25 : AO22x1_ASAP7_75t_R port map( A1 => header(14), A2 => granted_vc_1_port
                           , B1 => header(4), B2 => n7, Y => 
                           header_nxt_X_DEST_0_port);
   U26 : AO22x1_ASAP7_75t_R port map( A1 => header(19), A2 => granted_vc_1_port
                           , B1 => header(9), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_3_port);
   U27 : AO22x1_ASAP7_75t_R port map( A1 => header(18), A2 => granted_vc_1_port
                           , B1 => header(8), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_2_port);
   U28 : AO22x1_ASAP7_75t_R port map( A1 => header(17), A2 => granted_vc_1_port
                           , B1 => header(7), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_1_port);
   U29 : AO22x1_ASAP7_75t_R port map( A1 => header(16), A2 => granted_vc_1_port
                           , B1 => header(6), B2 => n7, Y => 
                           header_nxt_PACKET_LENGTH_0_port);
   rr_arbiter_no_delay_1 : rr_arbiter_no_delay_CNT2_6 port map( clk => clk, rst
                           => rst, req(1) => new_package_vc_1_port, req(0) => 
                           new_package_vc_0_port, ack => ack_vc, grant(1) => 
                           n13, grant(0) => granted_vc_0_port);
   routing_calc_1 : routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_6 port map( 
                           address(5) => header_nxt_X_DEST_1_port, address(4) 
                           => header_nxt_X_DEST_0_port, address(3) => 
                           header_nxt_Y_DEST_1_port, address(2) => 
                           header_nxt_Y_DEST_0_port, address(1) => 
                           header_nxt_Z_DEST_1_port, address(0) => 
                           header_nxt_Z_DEST_0_port, enable => routing_en, 
                           routing(6) => n_1502, routing(5) => 
                           granted_rq_5_port, routing(4) => n_1503, routing(3) 
                           => granted_rq_3, routing(2) => n_1504, routing(1) =>
                           n_1505, routing(0) => granted_rq_0);
   seq_packet_counter_i_0 : seq_packet_counter_1_12 port map( clk => clk, rst 
                           => rst, allocated => allocated_0_port, packet_len(3)
                           => header_nxt_PACKET_LENGTH_3_port, packet_len(2) =>
                           header_nxt_PACKET_LENGTH_2_port, packet_len(1) => 
                           header_nxt_PACKET_LENGTH_1_port, packet_len(0) => 
                           header_nxt_PACKET_LENGTH_0_port, enr_vc => enr_vc(0)
                           , flit_count(3) => flit_count_values_0_3_port, 
                           flit_count(2) => flit_count_values_0_2_port, 
                           flit_count(1) => flit_count_values_0_1_port, 
                           flit_count(0) => flit_count_values_0_0_port);
   seq_packet_counter_i_1 : seq_packet_counter_1_11 port map( clk => clk, rst 
                           => rst, allocated => allocated_1_port, packet_len(3)
                           => header_nxt_PACKET_LENGTH_3_port, packet_len(2) =>
                           header_nxt_PACKET_LENGTH_2_port, packet_len(1) => 
                           header_nxt_PACKET_LENGTH_1_port, packet_len(0) => 
                           header_nxt_PACKET_LENGTH_0_port, enr_vc => enr_vc(1)
                           , flit_count(3) => flit_count_values_1_3_port, 
                           flit_count(2) => flit_count_values_1_2_port, 
                           flit_count(1) => flit_count_values_1_1_port, 
                           flit_count(0) => flit_count_values_1_0_port);
   U3 : INVx1_ASAP7_75t_R port map( A => enr_vc(1), Y => n2);
   U4 : INVx1_ASAP7_75t_R port map( A => granted_vc_1_port, Y => n7);
   U5 : NOR2xp33_ASAP7_75t_R port map( A => n3, B => n8, Y => allocated_0_port)
                           ;
   U6 : NOR2xp33_ASAP7_75t_R port map( A => n7, B => n3, Y => allocated_1_port)
                           ;
   U7 : HB1xp67_ASAP7_75t_R port map( A => n13, Y => granted_vc_1_port);
   U8 : NOR4xp25_ASAP7_75t_R port map( A => flit_count_values_1_0_port, B => 
                           flit_count_values_1_1_port, C => 
                           flit_count_values_1_2_port, D => 
                           flit_count_values_1_3_port, Y => n10);
   U9 : NOR4xp25_ASAP7_75t_R port map( A => flit_count_values_0_0_port, B => 
                           flit_count_values_0_1_port, C => 
                           flit_count_values_0_2_port, D => 
                           flit_count_values_0_3_port, Y => n11);
   U10 : TIELOx1_ASAP7_75t_R port map( L => X_Logic0_port);
   U11 : INVx1_ASAP7_75t_R port map( A => ack_vc, Y => n3);
   U12 : INVx1_ASAP7_75t_R port map( A => enr_vc(0), Y => n4);
   U13 : INVx1_ASAP7_75t_R port map( A => flit_count_values_0_0_port, Y => n5);
   U14 : INVx1_ASAP7_75t_R port map( A => n11, Y => input_vc_in_use(0));
   U15 : INVx1_ASAP7_75t_R port map( A => granted_vc_0_port, Y => n8);
   U30 : INVx1_ASAP7_75t_R port map( A => flit_count_values_1_0_port, Y => n9);
   U31 : INVx1_ASAP7_75t_R port map( A => n10, Y => input_vc_in_use(1));

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity vc_output_allocator_port_num7_vc_num_out1 is

   port( clk, rst : in std_logic;  rq_vc_out : in std_logic_vector (5 downto 0)
         ;  granted_vc, packet_end : in std_logic_vector (11 downto 0);  
         crossbar_ctrl_vec : out std_logic_vector (2 downto 0);  vc_sel_enc, 
         output_vc_in_use : out std_logic;  ack_rq_vc_out : out 
         std_logic_vector (5 downto 0));

end vc_output_allocator_port_num7_vc_num_out1;

architecture SYN_rtl of vc_output_allocator_port_num7_vc_num_out1 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component rr_arbiter_no_delay_CNT6_0
      port( clk, rst : in std_logic;  req : in std_logic_vector (5 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (5 downto 0));
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI31xp33_ASAP7_75t_R
      port( A1, A2, A3, B : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1O1Ixp25_ASAP7_75t_R
      port( A1, A2, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal crossbar_ctrl_vec_2_port, crossbar_ctrl_vec_1_port, 
      crossbar_ctrl_vec_0_port, vc_sel_enc_0_0_port, output_vc_in_use_0_port, 
      grant_5_port, grant_4_port, grant_3_port, grant_2_port, grant_1_port, 
      grant_0_port, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18 : std_logic;

begin
   crossbar_ctrl_vec <= ( crossbar_ctrl_vec_2_port, crossbar_ctrl_vec_1_port, 
      crossbar_ctrl_vec_0_port );
   vc_sel_enc <= vc_sel_enc_0_0_port;
   output_vc_in_use <= output_vc_in_use_0_port;
   
   U13 : NAND2xp5_ASAP7_75t_R port map( A => vc_sel_enc_0_0_port, B => n25, Y 
                           => n26);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => n7, A2 => n2, B1 => n27, B2 => 
                           n25, Y => n51);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => n7, A2 => n16, B1 => n34, B2 => 
                           n25, Y => n52);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => n7, A2 => n17, B1 => n33, B2 => 
                           n25, Y => n53);
   U21 : NAND2xp5_ASAP7_75t_R port map( A => n14, B => n12, Y => n38);
   U22 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n39, A2 => n16, B => n40, C => 
                           n18, Y => n37);
   U23 : AOI22xp5_ASAP7_75t_R port map( A1 => packet_end(9), A2 => n2, B1 => 
                           packet_end(11), B2 => crossbar_ctrl_vec_0_port, Y =>
                           n39);
   U24 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n42, A2 => n16, B => n43, C => 
                           vc_sel_enc_0_0_port, Y => n36);
   U25 : AOI22xp5_ASAP7_75t_R port map( A1 => packet_end(8), A2 => n2, B1 => 
                           packet_end(10), B2 => crossbar_ctrl_vec_0_port, Y =>
                           n42);
   U26 : NAND2xp5_ASAP7_75t_R port map( A => n17, B => n16, Y => n47);
   U41 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n23, A2 => n24, B => n25, C =>
                           n26, Y => n50);
   U42 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(9), A2 => n27, B =>
                           n28, C => n11, Y => n24);
   U43 : AND2x2_ASAP7_75t_R port map( A => granted_vc(11), B => n10, Y => n28);
   U44 : A2O1A1O1Ixp25_ASAP7_75t_R port map( A1 => granted_vc(7), A2 => n10, B 
                           => n29, C => n13, D => n30, Y => n23);
   U45 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => granted_vc(1), A2 => n27, B =>
                           n32, C => n33, Y => n31);
   U46 : AND2x2_ASAP7_75t_R port map( A => granted_vc(3), B => n10, Y => n32);
   U47 : AND2x2_ASAP7_75t_R port map( A => granted_vc(5), B => n27, Y => n29);
   U48 : OAI31xp33_ASAP7_75t_R port map( A1 => n35, A2 => n36, A3 => n37, B => 
                           n25, Y => n54);
   U49 : OAI31xp33_ASAP7_75t_R port map( A1 => n38, A2 => grant_0_port, A3 => 
                           n10, B => n15, Y => n25);
   U50 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(5), A2 => n2, B => 
                           n41, C => crossbar_ctrl_vec_1_port, Y => n40);
   U51 : AND2x2_ASAP7_75t_R port map( A => packet_end(7), B => 
                           crossbar_ctrl_vec_0_port, Y => n41);
   U52 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(4), A2 => n2, B => 
                           n44, C => crossbar_ctrl_vec_1_port, Y => n43);
   U53 : AND2x2_ASAP7_75t_R port map( A => packet_end(6), B => 
                           crossbar_ctrl_vec_0_port, Y => n44);
   U54 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n45, A2 => n46, B => n47, C =>
                           output_vc_in_use_0_port, Y => n35);
   U55 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(0), A2 => n2, B => 
                           n48, C => n18, Y => n46);
   U56 : AND2x2_ASAP7_75t_R port map( A => packet_end(2), B => 
                           crossbar_ctrl_vec_0_port, Y => n48);
   U57 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => packet_end(1), A2 => n2, B => 
                           n49, C => vc_sel_enc_0_0_port, Y => n45);
   U58 : AND2x2_ASAP7_75t_R port map( A => packet_end(3), B => 
                           crossbar_ctrl_vec_0_port, Y => n49);
   U59 : AND2x2_ASAP7_75t_R port map( A => n15, B => grant_5_port, Y => 
                           ack_rq_vc_out(5));
   U60 : AND2x2_ASAP7_75t_R port map( A => n15, B => grant_3_port, Y => 
                           ack_rq_vc_out(3));
   U61 : AND2x2_ASAP7_75t_R port map( A => n15, B => grant_1_port, Y => 
                           ack_rq_vc_out(1));
   U62 : AND2x2_ASAP7_75t_R port map( A => n15, B => grant_0_port, Y => 
                           ack_rq_vc_out(0));
   rr_arbiter : rr_arbiter_no_delay_CNT6_0 port map( clk => clk, rst => rst, 
                           req(5) => rq_vc_out(5), req(4) => rq_vc_out(4), 
                           req(3) => rq_vc_out(3), req(2) => rq_vc_out(2), 
                           req(1) => rq_vc_out(1), req(0) => rq_vc_out(0), ack 
                           => n15, grant(5) => grant_5_port, grant(4) => 
                           grant_4_port, grant(3) => grant_3_port, grant(2) => 
                           grant_2_port, grant(1) => grant_1_port, grant(0) => 
                           grant_0_port);
   vc_sel_enc_int_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, 
                           CLK => clk, RESET => n3, SET => n1, QN => 
                           vc_sel_enc_0_0_port);
   crossbar_sels_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n5, CLK
                           => clk, RESET => n3, SET => n1, QN => 
                           crossbar_ctrl_vec_2_port);
   crossbar_sels_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n6, CLK
                           => clk, RESET => n3, SET => n1, QN => 
                           crossbar_ctrl_vec_1_port);
   crossbar_sels_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n4, CLK
                           => clk, RESET => n3, SET => n1, QN => 
                           crossbar_ctrl_vec_0_port);
   output_vc_in_use_int_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n9
                           , CLK => clk, RESET => n3, SET => n1, QN => 
                           output_vc_in_use_0_port);
   U3 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U4 : NOR2xp33_ASAP7_75t_R port map( A => n11, B => n31, Y => n30);
   U5 : NOR3xp33_ASAP7_75t_R port map( A => grant_3_port, B => grant_5_port, C 
                           => grant_1_port, Y => n27);
   U6 : NOR2xp33_ASAP7_75t_R port map( A => grant_5_port, B => grant_4_port, Y 
                           => n34);
   U7 : NOR2xp33_ASAP7_75t_R port map( A => grant_3_port, B => grant_2_port, Y 
                           => n33);
   U8 : INVx1_ASAP7_75t_R port map( A => rst, Y => n3);
   U9 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_0_port, Y => n2);
   U10 : NOR2xp33_ASAP7_75t_R port map( A => output_vc_in_use_0_port, B => n12,
                           Y => ack_rq_vc_out(4));
   U11 : NOR2xp33_ASAP7_75t_R port map( A => output_vc_in_use_0_port, B => n14,
                           Y => ack_rq_vc_out(2));
   U12 : INVx1_ASAP7_75t_R port map( A => n51, Y => n4);
   U14 : INVx1_ASAP7_75t_R port map( A => n52, Y => n5);
   U17 : INVx1_ASAP7_75t_R port map( A => n53, Y => n6);
   U19 : INVx1_ASAP7_75t_R port map( A => n25, Y => n7);
   U20 : INVx1_ASAP7_75t_R port map( A => n50, Y => n8);
   U27 : INVx1_ASAP7_75t_R port map( A => n54, Y => n9);
   U28 : INVx1_ASAP7_75t_R port map( A => n27, Y => n10);
   U29 : INVx1_ASAP7_75t_R port map( A => n34, Y => n11);
   U30 : INVx1_ASAP7_75t_R port map( A => grant_4_port, Y => n12);
   U31 : INVx1_ASAP7_75t_R port map( A => n33, Y => n13);
   U32 : INVx1_ASAP7_75t_R port map( A => grant_2_port, Y => n14);
   U33 : INVx1_ASAP7_75t_R port map( A => output_vc_in_use_0_port, Y => n15);
   U34 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_2_port, Y => n16);
   U35 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec_1_port, Y => n17);
   U36 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_0_0_port, Y => n18);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity header_arbiter_and_decoder_1_1_1_7_0_1_1_DXYU is

   port( clk, rst : in std_logic;  header : in std_logic_vector (9 downto 0);  
         valid_data_vc, enr_vc, ack_vc : in std_logic;  granted_rq : out 
         std_logic_vector (6 downto 0);  input_vc_in_use, packet_end, 
         granted_vc : out std_logic);

end header_arbiter_and_decoder_1_1_1_7_0_1_1_DXYU;

architecture SYN_rtl of header_arbiter_and_decoder_1_1_1_7_0_1_1_DXYU is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component NOR4xp25_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component seq_packet_counter_1_0
      port( clk, rst, allocated : in std_logic;  packet_len : in 
            std_logic_vector (3 downto 0);  enr_vc : in std_logic;  flit_count 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_0
      port( address : in std_logic_vector (5 downto 0);  enable : in std_logic;
            routing : out std_logic_vector (6 downto 0));
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR5xp2_ASAP7_75t_R
      port( A, B, C, D, E : in std_logic;  Y : out std_logic);
   end component;
   
   signal granted_vc_0_port, flit_count_values_0_3_port, 
      flit_count_values_0_2_port, flit_count_values_0_1_port, 
      flit_count_values_0_0_port, allocated_0_port, n4, n1, n2, n_1506 : 
      std_logic;

begin
   granted_vc <= granted_vc_0_port;
   
   U6 : NOR5xp2_ASAP7_75t_R port map( A => flit_count_values_0_2_port, B => 
                           flit_count_values_0_3_port, C => 
                           flit_count_values_0_1_port, D => n2, E => n1, Y => 
                           packet_end);
   U7 : AND2x2_ASAP7_75t_R port map( A => ack_vc, B => granted_vc_0_port, Y => 
                           allocated_0_port);
   U8 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc, B => n4, Y => 
                           granted_vc_0_port);
   routing_calc_1 : routing_calc_Xis1_Yis1_Zis1_rout_algoDXYU_0 port map( 
                           address(5) => header(5), address(4) => header(4), 
                           address(3) => header(3), address(2) => header(2), 
                           address(1) => header(1), address(0) => header(0), 
                           enable => granted_vc_0_port, routing(6) => 
                           granted_rq(6), routing(5) => granted_rq(5), 
                           routing(4) => granted_rq(4), routing(3) => 
                           granted_rq(3), routing(2) => granted_rq(2), 
                           routing(1) => granted_rq(1), routing(0) => n_1506);
   seq_packet_counter_i_0 : seq_packet_counter_1_0 port map( clk => clk, rst =>
                           rst, allocated => allocated_0_port, packet_len(3) =>
                           header(9), packet_len(2) => header(8), packet_len(1)
                           => header(7), packet_len(0) => header(6), enr_vc => 
                           enr_vc, flit_count(3) => flit_count_values_0_3_port,
                           flit_count(2) => flit_count_values_0_2_port, 
                           flit_count(1) => flit_count_values_0_1_port, 
                           flit_count(0) => flit_count_values_0_0_port);
   U2 : NOR4xp25_ASAP7_75t_R port map( A => flit_count_values_0_0_port, B => 
                           flit_count_values_0_1_port, C => 
                           flit_count_values_0_2_port, D => 
                           flit_count_values_0_3_port, Y => n4);
   U3 : TIELOx1_ASAP7_75t_R port map( L => granted_rq(0));
   U4 : INVx1_ASAP7_75t_R port map( A => enr_vc, Y => n1);
   U5 : INVx1_ASAP7_75t_R port map( A => flit_count_values_0_0_port, Y => n2);
   U9 : INVx1_ASAP7_75t_R port map( A => n4, Y => input_vc_in_use);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity switch_allocator_7_DXYU is

   port( clk, rst : in std_logic;  input_vc_in_use, output_vc_in_use : in 
         std_logic_vector (12 downto 0);  crossbar_ctrl_vec : in 
         std_logic_vector (38 downto 0);  vc_sel_enc_vec, valid_data_vc_vec, 
         incr_rx_vec : in std_logic_vector (12 downto 0);  crossbar_ctrl : out 
         std_logic_vector (20 downto 0);  vc_transfer_vec, vc_write_tx_vec : 
         out std_logic_vector (12 downto 0));

end switch_allocator_7_DXYU;

architecture SYN_rtl of switch_allocator_7_DXYU is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component TIEHIx1_ASAP7_75t_R
      port( H : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI31xp33_ASAP7_75t_R
      port( A1, A2, A3, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component HAxp5_ASAP7_75t_R
      port( A, B : in std_logic;  CON, SN : out std_logic);
   end component;
   
   component switch_allocator_7_DXYU_DW_mod_tc_6
      port( a : in std_logic_vector (4 downto 0);  b : in std_logic_vector (31 
            downto 0);  quotient : out std_logic_vector (4 downto 0);  
            remainder : out std_logic_vector (31 downto 0);  divide_by_0 : out 
            std_logic);
   end component;
   
   component switch_allocator_7_DXYU_DW_mod_tc_5
      port( a : in std_logic_vector (5 downto 0);  b : in std_logic_vector (31 
            downto 0);  quotient : out std_logic_vector (5 downto 0);  
            remainder : out std_logic_vector (31 downto 0);  divide_by_0 : out 
            std_logic);
   end component;
   
   component switch_allocator_7_DXYU_DW_mod_tc_4
      port( a : in std_logic_vector (5 downto 0);  b : in std_logic_vector (31 
            downto 0);  quotient : out std_logic_vector (5 downto 0);  
            remainder : out std_logic_vector (31 downto 0);  divide_by_0 : out 
            std_logic);
   end component;
   
   component switch_allocator_7_DXYU_DW_mod_tc_3
      port( a : in std_logic_vector (5 downto 0);  b : in std_logic_vector (31 
            downto 0);  quotient : out std_logic_vector (5 downto 0);  
            remainder : out std_logic_vector (31 downto 0);  divide_by_0 : out 
            std_logic);
   end component;
   
   component switch_allocator_7_DXYU_DW_mod_tc_2
      port( a : in std_logic_vector (5 downto 0);  b : in std_logic_vector (31 
            downto 0);  quotient : out std_logic_vector (5 downto 0);  
            remainder : out std_logic_vector (31 downto 0);  divide_by_0 : out 
            std_logic);
   end component;
   
   component switch_allocator_7_DXYU_DW_mod_tc_1
      port( a : in std_logic_vector (5 downto 0);  b : in std_logic_vector (31 
            downto 0);  quotient : out std_logic_vector (5 downto 0);  
            remainder : out std_logic_vector (31 downto 0);  divide_by_0 : out 
            std_logic);
   end component;
   
   component switch_allocator_7_DXYU_DW_mod_tc_0
      port( a : in std_logic_vector (5 downto 0);  b : in std_logic_vector (31 
            downto 0);  quotient : out std_logic_vector (5 downto 0);  
            remainder : out std_logic_vector (31 downto 0);  divide_by_0 : out 
            std_logic);
   end component;
   
   component credit_count_single_vc_depth_out2_1
      port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
            std_logic);
   end component;
   
   component credit_count_single_vc_depth_out2_2
      port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
            std_logic);
   end component;
   
   component rr_arbiter_no_delay_CNT2_7
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component credit_count_single_vc_depth_out2_3
      port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
            std_logic);
   end component;
   
   component credit_count_single_vc_depth_out2_4
      port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
            std_logic);
   end component;
   
   component rr_arbiter_no_delay_CNT2_8
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component credit_count_single_vc_depth_out2_5
      port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
            std_logic);
   end component;
   
   component credit_count_single_vc_depth_out2_6
      port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
            std_logic);
   end component;
   
   component rr_arbiter_no_delay_CNT2_9
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component credit_count_single_vc_depth_out2_7
      port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
            std_logic);
   end component;
   
   component credit_count_single_vc_depth_out2_8
      port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
            std_logic);
   end component;
   
   component rr_arbiter_no_delay_CNT2_10
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component credit_count_single_vc_depth_out2_9
      port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
            std_logic);
   end component;
   
   component credit_count_single_vc_depth_out2_10
      port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
            std_logic);
   end component;
   
   component rr_arbiter_no_delay_CNT2_11
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component credit_count_single_vc_depth_out2_11
      port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
            std_logic);
   end component;
   
   component credit_count_single_vc_depth_out2_12
      port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
            std_logic);
   end component;
   
   component rr_arbiter_no_delay_CNT2_12
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component credit_count_single_vc_depth_out2_0
      port( clk, rst, incr_rx, vc_write_tx : in std_logic;  credit_avail : out 
            std_logic);
   end component;
   
   component rr_arbiter_no_delay_CNT2_13
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component rr_arbiter_no_delay_CNT2_14
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component rr_arbiter_no_delay_CNT2_15
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component rr_arbiter_no_delay_CNT2_16
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component rr_arbiter_no_delay_CNT2_17
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component rr_arbiter_no_delay_CNT2_0
      port( clk, rst : in std_logic;  req : in std_logic_vector (1 downto 0);  
            ack : in std_logic;  grant : out std_logic_vector (1 downto 0));
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1O1Ixp25_ASAP7_75t_R
      port( A1, A2, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component A2O1A1Ixp33_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI322xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, B2, C1, C2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AND3x1_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OA211x2_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI32xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI33xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI333xp33_ASAP7_75t_R
      port( A1, A2, A3, B1, B2, B3, C1, C2, C3 : in std_logic;  Y : out 
            std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal n7, crossbar_ctrl_20_port, crossbar_ctrl_19_port, 
      crossbar_ctrl_18_port, crossbar_ctrl_17_port, crossbar_ctrl_16_port, 
      crossbar_ctrl_14_port, crossbar_ctrl_13_port, crossbar_ctrl_12_port, 
      crossbar_ctrl_8_port, crossbar_ctrl_7_port, crossbar_ctrl_6_port, 
      crossbar_ctrl_5_port, crossbar_ctrl_4_port, vc_write_tx_vec_12_port, 
      vc_write_tx_vec_11_port, vc_write_tx_vec_10_port, vc_write_tx_vec_9_port,
      vc_write_tx_vec_8_port, vc_write_tx_vec_7_port, vc_write_tx_vec_6_port, 
      vc_write_tx_vec_5_port, vc_write_tx_vec_4_port, vc_write_tx_vec_3_port, 
      vc_write_tx_vec_2_port, vc_write_tx_vec_1_port, switch_rq_12_port, 
      switch_rq_11_port, switch_rq_10_port, switch_rq_9_port, switch_rq_8_port,
      switch_rq_7_port, switch_rq_6_port, switch_rq_5_port, switch_rq_4_port, 
      switch_rq_3_port, switch_rq_2_port, switch_rq_1_port, 
      poss_channel_rq_6_5_1_port, poss_channel_rq_6_5_0_port, 
      poss_channel_rq_5_5_1_port, poss_channel_rq_5_5_0_port, 
      poss_channel_rq_5_4_1_port, poss_channel_rq_5_4_0_port, 
      poss_channel_rq_5_3_1_port, poss_channel_rq_5_3_0_port, 
      poss_channel_rq_5_2_1_port, poss_channel_rq_5_2_0_port, 
      poss_channel_rq_5_0_1_port, poss_channel_rq_5_0_0_port, 
      credit_avail_12_port, credit_avail_11_port, credit_avail_10_port, 
      credit_avail_9_port, credit_avail_8_port, credit_avail_7_port, 
      credit_avail_6_port, credit_avail_5_port, credit_avail_4_port, 
      credit_avail_3_port, credit_avail_2_port, credit_avail_1_port, 
      credit_avail_0_port, channel_rq_12_port, channel_rq_11_port, 
      channel_rq_10_port, channel_rq_9_port, channel_rq_8_port, 
      channel_rq_7_port, channel_rq_6_port, channel_rq_5_port, 
      channel_rq_4_port, channel_rq_3_port, channel_rq_2_port, 
      channel_rq_1_port, N0, N1, N2, N32, N33, N34, N64, N65, N66, N96, N97, 
      N98, N128, N129, N130, N160, N161, N162, N192, N193, N194, 
      switch_ack_var_6_port, switch_ack_var_5_port, switch_ack_var_4_port, 
      switch_ack_var_3_port, switch_ack_var_2_port, switch_ack_var_1_port, N426
      , N425, N401, N380, N379, N378, N377, N353, N330, N329, N309, N308, N307,
      net35534, n94, n95, n96_port, n97_port, n98_port, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128_port, n129_port, n130_port, n131, n132, n133, n134, n135, n136
      , n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160_port, n161_port, n162_port, n163, n164, n165, n166, n167, n168, n169
      , n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
      n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192_port, 
      n193_port, n194_port, n195, n196, n197, n198, n199, n200, n201, n202, 
      n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
      n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
      n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
      n239, n1_port, n2_port, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32_port, n33_port, n34_port, n35, n36, n37, n38, n39, n40, 
      n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, 
      vc_write_tx_vec_0_port, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
      n64_port, n65_port, n66_port, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
      n90, n91, n92, n93, n240, n241, n242, n243, n244, n245, n246, n247, n248,
      n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n_1507, 
      n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, 
      n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, 
      n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, 
      n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, 
      n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, 
      n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, 
      n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, 
      n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, 
      n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, 
      n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, 
      n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, 
      n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, 
      n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, 
      n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, 
      n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, 
      n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, 
      n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, 
      n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, 
      n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, 
      n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, 
      n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, 
      n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, 
      n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, 
      n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, 
      n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, 
      n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, 
      n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, 
      n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757 : std_logic;

begin
   crossbar_ctrl <= ( crossbar_ctrl_20_port, crossbar_ctrl_19_port, 
      crossbar_ctrl_18_port, crossbar_ctrl_17_port, crossbar_ctrl_16_port, N425
      , crossbar_ctrl_14_port, crossbar_ctrl_13_port, crossbar_ctrl_12_port, 
      N380, N378, N377, crossbar_ctrl_8_port, crossbar_ctrl_7_port, 
      crossbar_ctrl_6_port, crossbar_ctrl_5_port, crossbar_ctrl_4_port, N329, 
      crossbar_ctrl_vec(2), crossbar_ctrl_vec(1), crossbar_ctrl_vec(0) );
   vc_write_tx_vec <= ( vc_write_tx_vec_12_port, vc_write_tx_vec_11_port, 
      vc_write_tx_vec_10_port, vc_write_tx_vec_9_port, vc_write_tx_vec_8_port, 
      vc_write_tx_vec_7_port, vc_write_tx_vec_6_port, vc_write_tx_vec_5_port, 
      vc_write_tx_vec_4_port, vc_write_tx_vec_3_port, vc_write_tx_vec_2_port, 
      vc_write_tx_vec_1_port, vc_write_tx_vec_0_port );
   
   U35 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n141, A2 => n142, B => n258, C 
                           => n143, Y => n140);
   U37 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(0), A2 => n59
                           , B => n147, C => vc_sel_enc_vec(0), Y => n146);
   U38 : NAND2xp5_ASAP7_75t_R port map( A => poss_channel_rq_5_3_0_port, B => 
                           crossbar_ctrl_vec(0), Y => n147);
   U40 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(0), A2 => n73
                           , B => n148, C => n256, Y => n142);
   U41 : NAND2xp5_ASAP7_75t_R port map( A => poss_channel_rq_5_0_0_port, B => 
                           crossbar_ctrl_vec(0), Y => n148);
   U42 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(0), A2 => n67
                           , B => n149, C => n257, Y => n141);
   U43 : NAND2xp5_ASAP7_75t_R port map( A => poss_channel_rq_5_5_0_port, B => 
                           crossbar_ctrl_vec(0), Y => n149);
   U48 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n69, A2 => n241, B => n158, C 
                           => n93, Y => n157);
   U49 : NAND2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_vec(28), B => 
                           poss_channel_rq_5_3_1_port, Y => n158);
   U51 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(27), A2 => 
                           n59, B => n163, C => n240, Y => n162_port);
   U52 : NAND2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_vec(27), B => 
                           poss_channel_rq_5_3_0_port, Y => n163);
   U55 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n63, A2 => n91, B => n166, C =>
                           vc_sel_enc_vec(8), Y => n165);
   U56 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n61, A2 => n91, B => n167, C =>
                           n92, Y => n164);
   U57 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n63, A2 => n88, B => n170, C =>
                           vc_sel_enc_vec(7), Y => n169);
   U58 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n61, A2 => n88, B => n171, C =>
                           n89, Y => n168);
   U59 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(18), A2 => 
                           n59, B => n179, C => n85, Y => n178);
   U60 : NAND2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_vec(18), B => 
                           poss_channel_rq_5_3_0_port, Y => n179);
   U64 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(15), A2 => 
                           n59, B => n189, C => n82, Y => n188);
   U65 : NAND2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_vec(15), B => 
                           poss_channel_rq_5_3_0_port, Y => n189);
   U69 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n73, A2 => n79, B => n194_port,
                           C => vc_sel_enc_vec(4), Y => n193_port);
   U70 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(14), A2 => n249
                           , B1 => crossbar_ctrl_vec(12), B2 => 
                           poss_channel_rq_5_5_0_port, Y => n194_port);
   U71 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n69, A2 => n78, B => n195, C =>
                           n80, Y => n192_port);
   U72 : NAND2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_vec(13), B => 
                           poss_channel_rq_6_5_1_port, Y => n195);
   U73 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n70, A2 => n76, B => n198, C =>
                           vc_sel_enc_vec(3), Y => n197);
   U74 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(11), A2 => n249
                           , B1 => crossbar_ctrl_vec(10), B2 => 
                           poss_channel_rq_6_5_0_port, Y => n198);
   U75 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n69, A2 => n76, B => n199, C =>
                           n77, Y => n196);
   U76 : NAND2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_vec(10), B => 
                           poss_channel_rq_6_5_1_port, Y => n199);
   U77 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(6), A2 => n70
                           , B => n207, C => n254, Y => n206);
   U78 : NAND2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_vec(6), B => 
                           poss_channel_rq_6_5_0_port, Y => n207);
   U82 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(3), A2 => n70
                           , B => n217, C => n251, Y => n216);
   U83 : NAND2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_vec(3), B => 
                           poss_channel_rq_6_5_0_port, Y => n217);
   U88 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n73, A2 => n248, B => n223, C 
                           => vc_sel_enc_vec(12), Y => n222);
   U89 : NAND2xp5_ASAP7_75t_R port map( A => n249, B => n248, Y => n223);
   U92 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n73, A2 => n246, B => n227, C 
                           => vc_sel_enc_vec(11), Y => n226);
   U93 : NAND2xp5_ASAP7_75t_R port map( A => n249, B => n246, Y => n227);
   U95 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n69, A2 => n244, B => n234, C 
                           => n242, Y => n233);
   U96 : NAND2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_vec(31), B => 
                           poss_channel_rq_5_3_1_port, Y => n234);
   U98 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(30), A2 => 
                           n59, B => n239, C => n243, Y => n238);
   U99 : NAND2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_vec(30), B => 
                           poss_channel_rq_5_3_0_port, Y => n239);
   U102 : NAND2xp5_ASAP7_75t_R port map( A => valid_data_vc_vec(0), B => 
                           input_vc_in_use(0), Y => n97_port);
   U103 : OAI22xp5_ASAP7_75t_R port map( A1 => n71, A2 => n248, B1 => 
                           vc_write_tx_vec_11_port, B2 => n246, Y => 
                           crossbar_ctrl_18_port);
   U104 : OAI22xp5_ASAP7_75t_R port map( A1 => n244, A2 => n53, B1 => 
                           vc_write_tx_vec_9_port, B2 => n241, Y => 
                           crossbar_ctrl_17_port);
   U105 : OAI22xp5_ASAP7_75t_R port map( A1 => n53, A2 => n243, B1 => 
                           vc_write_tx_vec_9_port, B2 => n240, Y => 
                           crossbar_ctrl_16_port);
   U106 : OAI22xp5_ASAP7_75t_R port map( A1 => n53, A2 => n242, B1 => 
                           vc_write_tx_vec_9_port, B2 => n93, Y => N425);
   U107 : OAI22xp5_ASAP7_75t_R port map( A1 => n91, A2 => n60, B1 => 
                           vc_write_tx_vec_7_port, B2 => n88, Y => 
                           crossbar_ctrl_14_port);
   U108 : OAI22xp5_ASAP7_75t_R port map( A1 => n60, A2 => n90, B1 => 
                           vc_write_tx_vec_7_port, B2 => n87, Y => 
                           crossbar_ctrl_13_port);
   U109 : OAI22xp5_ASAP7_75t_R port map( A1 => n55, A2 => n85, B1 => 
                           vc_write_tx_vec_5_port, B2 => n82, Y => N380);
   U110 : OAI22xp5_ASAP7_75t_R port map( A1 => n84, A2 => n55, B1 => 
                           vc_write_tx_vec_5_port, B2 => n81, Y => N377);
   U111 : OAI22xp5_ASAP7_75t_R port map( A1 => vc_write_tx_vec_3_port, A2 => 
                           n76, B1 => n68, B2 => n78, Y => crossbar_ctrl_6_port
                           );
   U112 : OAI22xp5_ASAP7_75t_R port map( A1 => n62, A2 => n254, B1 => 
                           vc_write_tx_vec_1_port, B2 => n251, Y => 
                           crossbar_ctrl_4_port);
   U113 : OAI22xp5_ASAP7_75t_R port map( A1 => n62, A2 => n253, B1 => 
                           vc_write_tx_vec_1_port, B2 => n250, Y => N329);
   U200 : AOI333xp33_ASAP7_75t_R port map( A1 => n42, A2 => n41, A3 => n98_port
                           , B1 => n36, B2 => n35, B3 => n99, C1 => n39, C2 => 
                           n38, C3 => n100, Y => n96_port);
   U201 : AOI33xp33_ASAP7_75t_R port map( A1 => n45, A2 => n44, A3 => n101, B1 
                           => n48, B2 => n47, B3 => n102, Y => n95);
   U202 : AOI33xp33_ASAP7_75t_R port map( A1 => n51, A2 => n50, A3 => n103, B1 
                           => n34_port, B2 => n30, B3 => n104, Y => n94);
   U203 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc_vec(9), B => 
                           input_vc_in_use(9), Y => switch_rq_9_port);
   U204 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc_vec(8), B => 
                           input_vc_in_use(8), Y => switch_rq_8_port);
   U205 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc_vec(7), B => 
                           input_vc_in_use(7), Y => switch_rq_7_port);
   U206 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc_vec(6), B => 
                           input_vc_in_use(6), Y => switch_rq_6_port);
   U207 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc_vec(5), B => 
                           input_vc_in_use(5), Y => switch_rq_5_port);
   U208 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc_vec(4), B => 
                           input_vc_in_use(4), Y => switch_rq_4_port);
   U209 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc_vec(3), B => 
                           input_vc_in_use(3), Y => switch_rq_3_port);
   U210 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc_vec(2), B => 
                           input_vc_in_use(2), Y => switch_rq_2_port);
   U211 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc_vec(1), B => 
                           input_vc_in_use(1), Y => switch_rq_1_port);
   U212 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc_vec(12), B => 
                           input_vc_in_use(12), Y => switch_rq_12_port);
   U213 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc_vec(11), B => 
                           input_vc_in_use(11), Y => switch_rq_11_port);
   U214 : AND2x2_ASAP7_75t_R port map( A => valid_data_vc_vec(10), B => 
                           input_vc_in_use(10), Y => switch_rq_10_port);
   U215 : NAND3xp33_ASAP7_75t_R port map( A => n105, B => n106, C => n107, Y =>
                           switch_ack_var_6_port);
   U216 : AOI333xp33_ASAP7_75t_R port map( A1 => n108, A2 => n42, A3 => N97, B1
                           => n109, B2 => n36, B3 => N33, C1 => n110, C2 => n39
                           , C3 => N65, Y => n107);
   U217 : AOI33xp33_ASAP7_75t_R port map( A1 => n111, A2 => n45, A3 => N129, B1
                           => n112, B2 => n48, B3 => N161, Y => n106);
   U218 : AOI33xp33_ASAP7_75t_R port map( A1 => n113, A2 => n51, A3 => N193, B1
                           => n114, B2 => n34_port, B3 => N1, Y => n105);
   U219 : NAND3xp33_ASAP7_75t_R port map( A => n115, B => n116, C => n117, Y =>
                           switch_ack_var_5_port);
   U220 : AOI333xp33_ASAP7_75t_R port map( A1 => n108, A2 => n41, A3 => N96, B1
                           => n109, B2 => n35, B3 => N32, C1 => n110, C2 => n38
                           , C3 => N64, Y => n117);
   U221 : AOI33xp33_ASAP7_75t_R port map( A1 => n111, A2 => n44, A3 => N128, B1
                           => n112, B2 => n47, B3 => N160, Y => n116);
   U222 : AOI33xp33_ASAP7_75t_R port map( A1 => n113, A2 => n50, A3 => N192, B1
                           => n114, B2 => n30, B3 => N0, Y => n115);
   U223 : NAND3xp33_ASAP7_75t_R port map( A => n118, B => n119, C => n120, Y =>
                           switch_ack_var_4_port);
   U224 : AOI333xp33_ASAP7_75t_R port map( A1 => n42, A2 => n41, A3 => n108, B1
                           => n36, B2 => n35, B3 => n109, C1 => n39, C2 => n38,
                           C3 => n110, Y => n120);
   U225 : AOI33xp33_ASAP7_75t_R port map( A1 => n45, A2 => n44, A3 => n111, B1 
                           => n48, B2 => n47, B3 => n112, Y => n119);
   U226 : AOI33xp33_ASAP7_75t_R port map( A1 => n51, A2 => n50, A3 => n113, B1 
                           => n34_port, B2 => n30, B3 => n114, Y => n118);
   U227 : AND2x2_ASAP7_75t_R port map( A => N2, B => vc_write_tx_vec_0_port, Y 
                           => n114);
   U228 : NAND3xp33_ASAP7_75t_R port map( A => n128_port, B => n129_port, C => 
                           n130_port, Y => switch_ack_var_3_port);
   U229 : AOI333xp33_ASAP7_75t_R port map( A1 => n98_port, A2 => N96, A3 => N97
                           , B1 => n99, B2 => N32, B3 => N33, C1 => n100, C2 =>
                           N64, C3 => N65, Y => n130_port);
   U230 : AOI33xp33_ASAP7_75t_R port map( A1 => n101, A2 => N128, A3 => N129, 
                           B1 => n102, B2 => N160, B3 => N161, Y => n129_port);
   U231 : AOI33xp33_ASAP7_75t_R port map( A1 => n103, A2 => N192, A3 => N193, 
                           B1 => n104, B2 => N0, B3 => N1, Y => n128_port);
   U232 : NAND3xp33_ASAP7_75t_R port map( A => n131, B => n132, C => n133, Y =>
                           switch_ack_var_2_port);
   U233 : AOI333xp33_ASAP7_75t_R port map( A1 => n98_port, A2 => n42, A3 => N97
                           , B1 => n99, B2 => n36, B3 => N33, C1 => n100, C2 =>
                           n39, C3 => N65, Y => n133);
   U234 : AOI33xp33_ASAP7_75t_R port map( A1 => n101, A2 => n45, A3 => N129, B1
                           => n102, B2 => n48, B3 => N161, Y => n132);
   U235 : AOI33xp33_ASAP7_75t_R port map( A1 => n103, A2 => n51, A3 => N193, B1
                           => n104, B2 => n34_port, B3 => N1, Y => n131);
   U236 : NAND3xp33_ASAP7_75t_R port map( A => n134, B => n135, C => n136, Y =>
                           switch_ack_var_1_port);
   U237 : AOI333xp33_ASAP7_75t_R port map( A1 => N96, A2 => n41, A3 => n98_port
                           , B1 => N32, B2 => n35, B3 => n99, C1 => N64, C2 => 
                           n38, C3 => n100, Y => n136);
   U238 : AOI33xp33_ASAP7_75t_R port map( A1 => N128, A2 => n44, A3 => n101, B1
                           => N160, B2 => n47, B3 => n102, Y => n135);
   U239 : AOI33xp33_ASAP7_75t_R port map( A1 => N192, A2 => n50, A3 => n103, B1
                           => N0, B2 => n30, B3 => n104, Y => n134);
   U240 : NAND3xp33_ASAP7_75t_R port map( A => credit_avail_0_port, B => n137, 
                           C => output_vc_in_use(0), Y => n126);
   U241 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n138, A2 => n139, B => n258, 
                           C => n140, Y => n137);
   U242 : A2O1A1O1Ixp25_ASAP7_75t_R port map( A1 => poss_channel_rq_5_3_1_port,
                           A2 => crossbar_ctrl_vec(0), B => n145, C => 
                           vc_sel_enc_vec(0), D => n146, Y => n144);
   U243 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => poss_channel_rq_5_5_1_port, 
                           A2 => crossbar_ctrl_vec(0), B => n150, C => 
                           crossbar_ctrl_vec(1), Y => n139);
   U244 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => poss_channel_rq_5_0_1_port, 
                           A2 => crossbar_ctrl_vec(0), B => n151, C => 
                           crossbar_ctrl_vec(2), Y => n138);
   U245 : AND3x1_ASAP7_75t_R port map( A => credit_avail_9_port, B => n152, C 
                           => output_vc_in_use(9), Y => channel_rq_9_port);
   U246 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n153, A2 => n154, B => 
                           vc_sel_enc_vec(9), C => n155, Y => n152);
   U247 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n156, A2 => n93, B => n157, C
                           => vc_sel_enc_vec(9), Y => n155);
   U248 : OAI322xp33_ASAP7_75t_R port map( A1 => n74, A2 => 
                           crossbar_ctrl_vec(29), A3 => crossbar_ctrl_vec(28), 
                           B1 => n56, B2 => n240, C1 => n66_port, C2 => n241, Y
                           => n156);
   U249 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(27), A2 => 
                           poss_channel_rq_5_5_0_port, B => n159, C => 
                           crossbar_ctrl_vec(29), Y => n154);
   U250 : A2O1A1O1Ixp25_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(27), A2 
                           => n249, B => n160_port, C => n161_port, D => 
                           n162_port, Y => n153);
   U251 : OA211x2_ASAP7_75t_R port map( A1 => n164, A2 => n165, B => 
                           credit_avail_8_port, C => output_vc_in_use(8), Y => 
                           channel_rq_8_port);
   U252 : AOI32xp33_ASAP7_75t_R port map( A1 => n90, A2 => n91, A3 => 
                           poss_channel_rq_6_5_0_port, B1 => 
                           crossbar_ctrl_vec(25), B2 => n249, Y => n166);
   U253 : NAND3xp33_ASAP7_75t_R port map( A => n90, B => n91, C => 
                           poss_channel_rq_6_5_1_port, Y => n167);
   U254 : OA211x2_ASAP7_75t_R port map( A1 => n168, A2 => n169, B => 
                           credit_avail_7_port, C => output_vc_in_use(7), Y => 
                           channel_rq_7_port);
   U255 : AOI32xp33_ASAP7_75t_R port map( A1 => n87, A2 => n88, A3 => 
                           poss_channel_rq_6_5_0_port, B1 => 
                           crossbar_ctrl_vec(22), B2 => n249, Y => n170);
   U256 : NAND3xp33_ASAP7_75t_R port map( A => n87, B => n88, C => 
                           poss_channel_rq_6_5_1_port, Y => n171);
   U257 : AND3x1_ASAP7_75t_R port map( A => credit_avail_6_port, B => n172, C 
                           => output_vc_in_use(6), Y => channel_rq_6_port);
   U258 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n173, A2 => n174, B => n86, C
                           => n175, Y => n172);
   U259 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(19), A2 => 
                           n249, B => n57, C => n86, Y => n175);
   U260 : A2O1A1O1Ixp25_ASAP7_75t_R port map( A1 => poss_channel_rq_5_5_0_port,
                           A2 => n84, B => n177, C => n85, D => n178, Y => n176
                           );
   U261 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => poss_channel_rq_5_5_1_port, 
                           A2 => n84, B => n180, C => n85, Y => n174);
   U262 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(18), A2 => 
                           poss_channel_rq_5_3_1_port, B => n181, C => 
                           crossbar_ctrl_vec(20), Y => n173);
   U263 : AND3x1_ASAP7_75t_R port map( A => credit_avail_5_port, B => n182, C 
                           => output_vc_in_use(5), Y => channel_rq_5_port);
   U264 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n183, A2 => n184, B => n83, C
                           => n185, Y => n182);
   U265 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(16), A2 => 
                           n249, B => n58, C => n83, Y => n185);
   U266 : A2O1A1O1Ixp25_ASAP7_75t_R port map( A1 => poss_channel_rq_5_5_0_port,
                           A2 => n81, B => n187, C => n82, D => n188, Y => n186
                           );
   U267 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => poss_channel_rq_5_5_1_port, 
                           A2 => n81, B => n190, C => n82, Y => n184);
   U268 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(15), A2 => 
                           poss_channel_rq_5_3_1_port, B => n191, C => 
                           crossbar_ctrl_vec(17), Y => n183);
   U269 : OA211x2_ASAP7_75t_R port map( A1 => n192_port, A2 => n193_port, B => 
                           credit_avail_4_port, C => output_vc_in_use(4), Y => 
                           channel_rq_4_port);
   U270 : OA211x2_ASAP7_75t_R port map( A1 => n196, A2 => n197, B => 
                           credit_avail_3_port, C => output_vc_in_use(3), Y => 
                           channel_rq_3_port);
   U271 : AND3x1_ASAP7_75t_R port map( A => credit_avail_2_port, B => n200, C 
                           => output_vc_in_use(2), Y => channel_rq_2_port);
   U272 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n201, A2 => n202, B => n255, 
                           C => n203, Y => n200);
   U273 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(8), A2 => 
                           n249, B => n64_port, C => n255, Y => n203);
   U274 : A2O1A1O1Ixp25_ASAP7_75t_R port map( A1 => poss_channel_rq_5_3_0_port,
                           A2 => n253, B => n205, C => n254, D => n206, Y => 
                           n204);
   U275 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => poss_channel_rq_5_3_1_port, 
                           A2 => n253, B => n208, C => n254, Y => n202);
   U276 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(6), A2 => 
                           poss_channel_rq_6_5_1_port, B => n209, C => 
                           crossbar_ctrl_vec(7), Y => n201);
   U277 : AND3x1_ASAP7_75t_R port map( A => credit_avail_1_port, B => n210, C 
                           => output_vc_in_use(1), Y => channel_rq_1_port);
   U278 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n211, A2 => n212, B => n252, 
                           C => n213, Y => n210);
   U279 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(5), A2 => 
                           n249, B => n65_port, C => n252, Y => n213);
   U280 : A2O1A1O1Ixp25_ASAP7_75t_R port map( A1 => poss_channel_rq_5_3_0_port,
                           A2 => n250, B => n215, C => n251, D => n216, Y => 
                           n214);
   U281 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => poss_channel_rq_5_3_1_port, 
                           A2 => n250, B => n218, C => n251, Y => n212);
   U282 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(3), A2 => 
                           poss_channel_rq_6_5_1_port, B => n219, C => 
                           crossbar_ctrl_vec(4), Y => n211);
   U283 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n221, A2 => 
                           vc_sel_enc_vec(12), B => n222, C => 
                           credit_avail_12_port, Y => n220);
   U284 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n225, A2 => 
                           vc_sel_enc_vec(11), B => n226, C => 
                           credit_avail_11_port, Y => n224);
   U285 : AND3x1_ASAP7_75t_R port map( A => credit_avail_10_port, B => n228, C 
                           => output_vc_in_use(10), Y => channel_rq_10_port);
   U286 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n229, A2 => n230, B => 
                           vc_sel_enc_vec(10), C => n231, Y => n228);
   U287 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => n232, A2 => n242, B => n233, 
                           C => vc_sel_enc_vec(10), Y => n231);
   U288 : OAI322xp33_ASAP7_75t_R port map( A1 => n74, A2 => 
                           crossbar_ctrl_vec(32), A3 => crossbar_ctrl_vec(31), 
                           B1 => n56, B2 => n243, C1 => n66_port, C2 => n244, Y
                           => n232);
   U289 : A2O1A1Ixp33_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(30), A2 => 
                           poss_channel_rq_5_5_0_port, B => n235, C => 
                           crossbar_ctrl_vec(32), Y => n230);
   U290 : A2O1A1O1Ixp25_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(30), A2 
                           => n249, B => n236, C => n237, D => n238, Y => n229)
                           ;
   U291 : AO22x1_ASAP7_75t_R port map( A1 => vc_write_tx_vec_11_port, A2 => 
                           crossbar_ctrl_vec(38), B1 => crossbar_ctrl_vec(35), 
                           B2 => n71, Y => crossbar_ctrl_20_port);
   U292 : AO22x1_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(37), A2 => 
                           vc_write_tx_vec_11_port, B1 => crossbar_ctrl_vec(34)
                           , B2 => n71, Y => crossbar_ctrl_19_port);
   U293 : AO22x1_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(24), A2 => 
                           vc_write_tx_vec_7_port, B1 => crossbar_ctrl_vec(21),
                           B2 => n60, Y => crossbar_ctrl_12_port);
   U294 : AO22x1_ASAP7_75t_R port map( A1 => vc_write_tx_vec_5_port, A2 => 
                           crossbar_ctrl_vec(19), B1 => n55, B2 => 
                           crossbar_ctrl_vec(16), Y => N378);
   U295 : AO22x1_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(14), A2 => 
                           vc_write_tx_vec_3_port, B1 => n68, B2 => 
                           crossbar_ctrl_vec(11), Y => crossbar_ctrl_8_port);
   U296 : AO22x1_ASAP7_75t_R port map( A1 => vc_write_tx_vec_3_port, A2 => 
                           crossbar_ctrl_vec(13), B1 => n68, B2 => 
                           crossbar_ctrl_vec(10), Y => crossbar_ctrl_7_port);
   U297 : AO22x1_ASAP7_75t_R port map( A1 => crossbar_ctrl_vec(8), A2 => 
                           vc_write_tx_vec_1_port, B1 => n62, B2 => 
                           crossbar_ctrl_vec(5), Y => crossbar_ctrl_5_port);
   rr_arbiter_1 : rr_arbiter_no_delay_CNT2_0 port map( clk => clk, rst => rst, 
                           req(1) => switch_rq_2_port, req(0) => 
                           switch_rq_1_port, ack => switch_ack_var_1_port, 
                           grant(1) => poss_channel_rq_5_2_1_port, grant(0) => 
                           poss_channel_rq_5_2_0_port);
   rr_arbiter_2 : rr_arbiter_no_delay_CNT2_17 port map( clk => clk, rst => n21,
                           req(1) => switch_rq_4_port, req(0) => 
                           switch_rq_3_port, ack => switch_ack_var_2_port, 
                           grant(1) => poss_channel_rq_5_3_1_port, grant(0) => 
                           poss_channel_rq_5_3_0_port);
   rr_arbiter_3 : rr_arbiter_no_delay_CNT2_16 port map( clk => clk, rst => n21,
                           req(1) => switch_rq_6_port, req(0) => 
                           switch_rq_5_port, ack => switch_ack_var_3_port, 
                           grant(1) => poss_channel_rq_5_4_1_port, grant(0) => 
                           poss_channel_rq_5_4_0_port);
   rr_arbiter_4 : rr_arbiter_no_delay_CNT2_15 port map( clk => clk, rst => n21,
                           req(1) => switch_rq_8_port, req(0) => 
                           switch_rq_7_port, ack => switch_ack_var_4_port, 
                           grant(1) => poss_channel_rq_5_5_1_port, grant(0) => 
                           poss_channel_rq_5_5_0_port);
   rr_arbiter_5 : rr_arbiter_no_delay_CNT2_14 port map( clk => clk, rst => n21,
                           req(1) => switch_rq_10_port, req(0) => 
                           switch_rq_9_port, ack => switch_ack_var_5_port, 
                           grant(1) => poss_channel_rq_6_5_1_port, grant(0) => 
                           poss_channel_rq_6_5_0_port);
   rr_arbiter_6 : rr_arbiter_no_delay_CNT2_13 port map( clk => clk, rst => n21,
                           req(1) => switch_rq_12_port, req(0) => 
                           switch_rq_11_port, ack => switch_ack_var_6_port, 
                           grant(1) => poss_channel_rq_5_0_1_port, grant(0) => 
                           poss_channel_rq_5_0_0_port);
   credit_count_i_0_0 : credit_count_single_vc_depth_out2_0 port map( clk => 
                           clk, rst => n21, incr_rx => incr_rx_vec(0), 
                           vc_write_tx => vc_write_tx_vec_0_port, credit_avail 
                           => credit_avail_0_port);
   rr_arbiter_1_0 : rr_arbiter_no_delay_CNT2_12 port map( clk => clk, rst => 
                           n21, req(1) => channel_rq_2_port, req(0) => 
                           channel_rq_1_port, ack => n7, grant(1) => 
                           vc_write_tx_vec_2_port, grant(0) => 
                           vc_write_tx_vec_1_port);
   credit_count_i_1_1 : credit_count_single_vc_depth_out2_12 port map( clk => 
                           clk, rst => n20, incr_rx => incr_rx_vec(1), 
                           vc_write_tx => vc_write_tx_vec_1_port, credit_avail 
                           => credit_avail_1_port);
   credit_count_i_1_2 : credit_count_single_vc_depth_out2_11 port map( clk => 
                           clk, rst => n20, incr_rx => incr_rx_vec(2), 
                           vc_write_tx => vc_write_tx_vec_2_port, credit_avail 
                           => credit_avail_2_port);
   rr_arbiter_2_0 : rr_arbiter_no_delay_CNT2_11 port map( clk => clk, rst => 
                           n21, req(1) => channel_rq_4_port, req(0) => 
                           channel_rq_3_port, ack => n7, grant(1) => 
                           vc_write_tx_vec_4_port, grant(0) => 
                           vc_write_tx_vec_3_port);
   credit_count_i_2_3 : credit_count_single_vc_depth_out2_10 port map( clk => 
                           clk, rst => n20, incr_rx => incr_rx_vec(3), 
                           vc_write_tx => vc_write_tx_vec_3_port, credit_avail 
                           => credit_avail_3_port);
   credit_count_i_2_4 : credit_count_single_vc_depth_out2_9 port map( clk => 
                           clk, rst => n20, incr_rx => incr_rx_vec(4), 
                           vc_write_tx => vc_write_tx_vec_4_port, credit_avail 
                           => credit_avail_4_port);
   rr_arbiter_3_0 : rr_arbiter_no_delay_CNT2_10 port map( clk => clk, rst => 
                           n21, req(1) => channel_rq_6_port, req(0) => 
                           channel_rq_5_port, ack => n7, grant(1) => 
                           vc_write_tx_vec_6_port, grant(0) => 
                           vc_write_tx_vec_5_port);
   credit_count_i_3_5 : credit_count_single_vc_depth_out2_8 port map( clk => 
                           clk, rst => n20, incr_rx => incr_rx_vec(5), 
                           vc_write_tx => vc_write_tx_vec_5_port, credit_avail 
                           => credit_avail_5_port);
   credit_count_i_3_6 : credit_count_single_vc_depth_out2_7 port map( clk => 
                           clk, rst => n20, incr_rx => incr_rx_vec(6), 
                           vc_write_tx => vc_write_tx_vec_6_port, credit_avail 
                           => credit_avail_6_port);
   rr_arbiter_4_0 : rr_arbiter_no_delay_CNT2_9 port map( clk => clk, rst => n21
                           , req(1) => channel_rq_8_port, req(0) => 
                           channel_rq_7_port, ack => n7, grant(1) => 
                           vc_write_tx_vec_8_port, grant(0) => 
                           vc_write_tx_vec_7_port);
   credit_count_i_4_7 : credit_count_single_vc_depth_out2_6 port map( clk => 
                           clk, rst => n20, incr_rx => incr_rx_vec(7), 
                           vc_write_tx => vc_write_tx_vec_7_port, credit_avail 
                           => credit_avail_7_port);
   credit_count_i_4_8 : credit_count_single_vc_depth_out2_5 port map( clk => 
                           clk, rst => n20, incr_rx => incr_rx_vec(8), 
                           vc_write_tx => vc_write_tx_vec_8_port, credit_avail 
                           => credit_avail_8_port);
   rr_arbiter_5_0 : rr_arbiter_no_delay_CNT2_8 port map( clk => clk, rst => n21
                           , req(1) => channel_rq_10_port, req(0) => 
                           channel_rq_9_port, ack => n7, grant(1) => 
                           vc_write_tx_vec_10_port, grant(0) => 
                           vc_write_tx_vec_9_port);
   credit_count_i_5_9 : credit_count_single_vc_depth_out2_4 port map( clk => 
                           clk, rst => n20, incr_rx => incr_rx_vec(9), 
                           vc_write_tx => vc_write_tx_vec_9_port, credit_avail 
                           => credit_avail_9_port);
   credit_count_i_5_10 : credit_count_single_vc_depth_out2_3 port map( clk => 
                           clk, rst => n20, incr_rx => incr_rx_vec(10), 
                           vc_write_tx => vc_write_tx_vec_10_port, credit_avail
                           => credit_avail_10_port);
   rr_arbiter_6_0 : rr_arbiter_no_delay_CNT2_7 port map( clk => clk, rst => n21
                           , req(1) => channel_rq_12_port, req(0) => 
                           channel_rq_11_port, ack => n7, grant(1) => 
                           vc_write_tx_vec_12_port, grant(0) => 
                           vc_write_tx_vec_11_port);
   credit_count_i_6_11 : credit_count_single_vc_depth_out2_2 port map( clk => 
                           clk, rst => n20, incr_rx => incr_rx_vec(11), 
                           vc_write_tx => vc_write_tx_vec_11_port, credit_avail
                           => credit_avail_11_port);
   credit_count_i_6_12 : credit_count_single_vc_depth_out2_1 port map( clk => 
                           clk, rst => n20, incr_rx => incr_rx_vec(12), 
                           vc_write_tx => vc_write_tx_vec_12_port, credit_avail
                           => credit_avail_12_port);
   mod_219_G7 : switch_allocator_7_DXYU_DW_mod_tc_0 port map( a(5) => net35534,
                           a(4) => net35534, a(3) => n13, a(2) => n3, a(1) => 
                           n14, a(0) => n19, b(31) => net35534, b(30) => 
                           net35534, b(29) => net35534, b(28) => net35534, 
                           b(27) => net35534, b(26) => net35534, b(25) => 
                           net35534, b(24) => net35534, b(23) => net35534, 
                           b(22) => net35534, b(21) => net35534, b(20) => 
                           net35534, b(19) => net35534, b(18) => net35534, 
                           b(17) => net35534, b(16) => net35534, b(15) => 
                           net35534, b(14) => net35534, b(13) => net35534, 
                           b(12) => net35534, b(11) => net35534, b(10) => 
                           net35534, b(9) => net35534, b(8) => net35534, b(7) 
                           => net35534, b(6) => net35534, b(5) => net35534, 
                           b(4) => net35534, b(3) => net35534, b(2) => n7, b(1)
                           => n7, b(0) => n7, quotient(5) => n_1508, 
                           quotient(4) => n_1509, quotient(3) => n_1510, 
                           quotient(2) => n_1511, quotient(1) => n_1512, 
                           quotient(0) => n_1513, remainder(31) => n_1514, 
                           remainder(30) => n_1515, remainder(29) => n_1516, 
                           remainder(28) => n_1517, remainder(27) => n_1518, 
                           remainder(26) => n_1519, remainder(25) => n_1520, 
                           remainder(24) => n_1521, remainder(23) => n_1522, 
                           remainder(22) => n_1523, remainder(21) => n_1524, 
                           remainder(20) => n_1525, remainder(19) => n_1526, 
                           remainder(18) => n_1527, remainder(17) => n_1528, 
                           remainder(16) => n_1529, remainder(15) => n_1530, 
                           remainder(14) => n_1531, remainder(13) => n_1532, 
                           remainder(12) => n_1533, remainder(11) => n_1534, 
                           remainder(10) => n_1535, remainder(9) => n_1536, 
                           remainder(8) => n_1537, remainder(7) => n_1538, 
                           remainder(6) => n_1539, remainder(5) => n_1540, 
                           remainder(4) => n_1541, remainder(3) => n_1542, 
                           remainder(2) => N194, remainder(1) => N193, 
                           remainder(0) => N192, divide_by_0 => n_1507);
   mod_219_G6 : switch_allocator_7_DXYU_DW_mod_tc_1 port map( a(5) => net35534,
                           a(4) => net35534, a(3) => n16, a(2) => n11, a(1) => 
                           N426, a(0) => N425, b(31) => net35534, b(30) => 
                           net35534, b(29) => net35534, b(28) => net35534, 
                           b(27) => net35534, b(26) => net35534, b(25) => 
                           net35534, b(24) => net35534, b(23) => net35534, 
                           b(22) => net35534, b(21) => net35534, b(20) => 
                           net35534, b(19) => net35534, b(18) => net35534, 
                           b(17) => net35534, b(16) => net35534, b(15) => 
                           net35534, b(14) => net35534, b(13) => net35534, 
                           b(12) => net35534, b(11) => net35534, b(10) => 
                           net35534, b(9) => net35534, b(8) => net35534, b(7) 
                           => net35534, b(6) => net35534, b(5) => net35534, 
                           b(4) => net35534, b(3) => net35534, b(2) => n7, b(1)
                           => n7, b(0) => n7, quotient(5) => n_1544, 
                           quotient(4) => n_1545, quotient(3) => n_1546, 
                           quotient(2) => n_1547, quotient(1) => n_1548, 
                           quotient(0) => n_1549, remainder(31) => n_1550, 
                           remainder(30) => n_1551, remainder(29) => n_1552, 
                           remainder(28) => n_1553, remainder(27) => n_1554, 
                           remainder(26) => n_1555, remainder(25) => n_1556, 
                           remainder(24) => n_1557, remainder(23) => n_1558, 
                           remainder(22) => n_1559, remainder(21) => n_1560, 
                           remainder(20) => n_1561, remainder(19) => n_1562, 
                           remainder(18) => n_1563, remainder(17) => n_1564, 
                           remainder(16) => n_1565, remainder(15) => n_1566, 
                           remainder(14) => n_1567, remainder(13) => n_1568, 
                           remainder(12) => n_1569, remainder(11) => n_1570, 
                           remainder(10) => n_1571, remainder(9) => n_1572, 
                           remainder(8) => n_1573, remainder(7) => n_1574, 
                           remainder(6) => n_1575, remainder(5) => n_1576, 
                           remainder(4) => n_1577, remainder(3) => n_1578, 
                           remainder(2) => N162, remainder(1) => N161, 
                           remainder(0) => N160, divide_by_0 => n_1543);
   mod_219_G5 : switch_allocator_7_DXYU_DW_mod_tc_2 port map( a(5) => net35534,
                           a(4) => net35534, a(3) => n17, a(2) => n2_port, a(1)
                           => n15, a(0) => N401, b(31) => net35534, b(30) => 
                           net35534, b(29) => net35534, b(28) => net35534, 
                           b(27) => net35534, b(26) => net35534, b(25) => 
                           net35534, b(24) => net35534, b(23) => net35534, 
                           b(22) => net35534, b(21) => net35534, b(20) => 
                           net35534, b(19) => net35534, b(18) => net35534, 
                           b(17) => net35534, b(16) => net35534, b(15) => 
                           net35534, b(14) => net35534, b(13) => net35534, 
                           b(12) => net35534, b(11) => net35534, b(10) => 
                           net35534, b(9) => net35534, b(8) => net35534, b(7) 
                           => net35534, b(6) => net35534, b(5) => net35534, 
                           b(4) => net35534, b(3) => net35534, b(2) => n7, b(1)
                           => n7, b(0) => n7, quotient(5) => n_1580, 
                           quotient(4) => n_1581, quotient(3) => n_1582, 
                           quotient(2) => n_1583, quotient(1) => n_1584, 
                           quotient(0) => n_1585, remainder(31) => n_1586, 
                           remainder(30) => n_1587, remainder(29) => n_1588, 
                           remainder(28) => n_1589, remainder(27) => n_1590, 
                           remainder(26) => n_1591, remainder(25) => n_1592, 
                           remainder(24) => n_1593, remainder(23) => n_1594, 
                           remainder(22) => n_1595, remainder(21) => n_1596, 
                           remainder(20) => n_1597, remainder(19) => n_1598, 
                           remainder(18) => n_1599, remainder(17) => n_1600, 
                           remainder(16) => n_1601, remainder(15) => n_1602, 
                           remainder(14) => n_1603, remainder(13) => n_1604, 
                           remainder(12) => n_1605, remainder(11) => n_1606, 
                           remainder(10) => n_1607, remainder(9) => n_1608, 
                           remainder(8) => n_1609, remainder(7) => n_1610, 
                           remainder(6) => n_1611, remainder(5) => n_1612, 
                           remainder(4) => n_1613, remainder(3) => n_1614, 
                           remainder(2) => N130, remainder(1) => N129, 
                           remainder(0) => N128, divide_by_0 => n_1579);
   mod_219_G4 : switch_allocator_7_DXYU_DW_mod_tc_3 port map( a(5) => net35534,
                           a(4) => net35534, a(3) => N380, a(2) => N379, a(1) 
                           => N378, a(0) => N377, b(31) => net35534, b(30) => 
                           net35534, b(29) => net35534, b(28) => net35534, 
                           b(27) => net35534, b(26) => net35534, b(25) => 
                           net35534, b(24) => net35534, b(23) => net35534, 
                           b(22) => net35534, b(21) => net35534, b(20) => 
                           net35534, b(19) => net35534, b(18) => net35534, 
                           b(17) => net35534, b(16) => net35534, b(15) => 
                           net35534, b(14) => net35534, b(13) => net35534, 
                           b(12) => net35534, b(11) => net35534, b(10) => 
                           net35534, b(9) => net35534, b(8) => net35534, b(7) 
                           => net35534, b(6) => net35534, b(5) => net35534, 
                           b(4) => net35534, b(3) => net35534, b(2) => n7, b(1)
                           => n7, b(0) => n7, quotient(5) => n_1616, 
                           quotient(4) => n_1617, quotient(3) => n_1618, 
                           quotient(2) => n_1619, quotient(1) => n_1620, 
                           quotient(0) => n_1621, remainder(31) => n_1622, 
                           remainder(30) => n_1623, remainder(29) => n_1624, 
                           remainder(28) => n_1625, remainder(27) => n_1626, 
                           remainder(26) => n_1627, remainder(25) => n_1628, 
                           remainder(24) => n_1629, remainder(23) => n_1630, 
                           remainder(22) => n_1631, remainder(21) => n_1632, 
                           remainder(20) => n_1633, remainder(19) => n_1634, 
                           remainder(18) => n_1635, remainder(17) => n_1636, 
                           remainder(16) => n_1637, remainder(15) => n_1638, 
                           remainder(14) => n_1639, remainder(13) => n_1640, 
                           remainder(12) => n_1641, remainder(11) => n_1642, 
                           remainder(10) => n_1643, remainder(9) => n_1644, 
                           remainder(8) => n_1645, remainder(7) => n_1646, 
                           remainder(6) => n_1647, remainder(5) => n_1648, 
                           remainder(4) => n_1649, remainder(3) => n_1650, 
                           remainder(2) => N98, remainder(1) => N97, 
                           remainder(0) => N96, divide_by_0 => n_1615);
   mod_219_G3 : switch_allocator_7_DXYU_DW_mod_tc_4 port map( a(5) => net35534,
                           a(4) => net35534, a(3) => n10, a(2) => n1_port, a(1)
                           => n9, a(0) => N353, b(31) => net35534, b(30) => 
                           net35534, b(29) => net35534, b(28) => net35534, 
                           b(27) => net35534, b(26) => net35534, b(25) => 
                           net35534, b(24) => net35534, b(23) => net35534, 
                           b(22) => net35534, b(21) => net35534, b(20) => 
                           net35534, b(19) => net35534, b(18) => net35534, 
                           b(17) => net35534, b(16) => net35534, b(15) => 
                           net35534, b(14) => net35534, b(13) => net35534, 
                           b(12) => net35534, b(11) => net35534, b(10) => 
                           net35534, b(9) => net35534, b(8) => net35534, b(7) 
                           => net35534, b(6) => net35534, b(5) => net35534, 
                           b(4) => net35534, b(3) => net35534, b(2) => n7, b(1)
                           => n7, b(0) => n7, quotient(5) => n_1652, 
                           quotient(4) => n_1653, quotient(3) => n_1654, 
                           quotient(2) => n_1655, quotient(1) => n_1656, 
                           quotient(0) => n_1657, remainder(31) => n_1658, 
                           remainder(30) => n_1659, remainder(29) => n_1660, 
                           remainder(28) => n_1661, remainder(27) => n_1662, 
                           remainder(26) => n_1663, remainder(25) => n_1664, 
                           remainder(24) => n_1665, remainder(23) => n_1666, 
                           remainder(22) => n_1667, remainder(21) => n_1668, 
                           remainder(20) => n_1669, remainder(19) => n_1670, 
                           remainder(18) => n_1671, remainder(17) => n_1672, 
                           remainder(16) => n_1673, remainder(15) => n_1674, 
                           remainder(14) => n_1675, remainder(13) => n_1676, 
                           remainder(12) => n_1677, remainder(11) => n_1678, 
                           remainder(10) => n_1679, remainder(9) => n_1680, 
                           remainder(8) => n_1681, remainder(7) => n_1682, 
                           remainder(6) => n_1683, remainder(5) => n_1684, 
                           remainder(4) => n_1685, remainder(3) => n_1686, 
                           remainder(2) => N66, remainder(1) => N65, 
                           remainder(0) => N64, divide_by_0 => n_1651);
   mod_219_G2 : switch_allocator_7_DXYU_DW_mod_tc_5 port map( a(5) => net35534,
                           a(4) => net35534, a(3) => n12, a(2) => n5, a(1) => 
                           N330, a(0) => N329, b(31) => net35534, b(30) => 
                           net35534, b(29) => net35534, b(28) => net35534, 
                           b(27) => net35534, b(26) => net35534, b(25) => 
                           net35534, b(24) => net35534, b(23) => net35534, 
                           b(22) => net35534, b(21) => net35534, b(20) => 
                           net35534, b(19) => net35534, b(18) => net35534, 
                           b(17) => net35534, b(16) => net35534, b(15) => 
                           net35534, b(14) => net35534, b(13) => net35534, 
                           b(12) => net35534, b(11) => net35534, b(10) => 
                           net35534, b(9) => net35534, b(8) => net35534, b(7) 
                           => net35534, b(6) => net35534, b(5) => net35534, 
                           b(4) => net35534, b(3) => net35534, b(2) => n7, b(1)
                           => n7, b(0) => n7, quotient(5) => n_1688, 
                           quotient(4) => n_1689, quotient(3) => n_1690, 
                           quotient(2) => n_1691, quotient(1) => n_1692, 
                           quotient(0) => n_1693, remainder(31) => n_1694, 
                           remainder(30) => n_1695, remainder(29) => n_1696, 
                           remainder(28) => n_1697, remainder(27) => n_1698, 
                           remainder(26) => n_1699, remainder(25) => n_1700, 
                           remainder(24) => n_1701, remainder(23) => n_1702, 
                           remainder(22) => n_1703, remainder(21) => n_1704, 
                           remainder(20) => n_1705, remainder(19) => n_1706, 
                           remainder(18) => n_1707, remainder(17) => n_1708, 
                           remainder(16) => n_1709, remainder(15) => n_1710, 
                           remainder(14) => n_1711, remainder(13) => n_1712, 
                           remainder(12) => n_1713, remainder(11) => n_1714, 
                           remainder(10) => n_1715, remainder(9) => n_1716, 
                           remainder(8) => n_1717, remainder(7) => n_1718, 
                           remainder(6) => n_1719, remainder(5) => n_1720, 
                           remainder(4) => n_1721, remainder(3) => n_1722, 
                           remainder(2) => N34, remainder(1) => N33, 
                           remainder(0) => N32, divide_by_0 => n_1687);
   mod_219 : switch_allocator_7_DXYU_DW_mod_tc_6 port map( a(4) => net35534, 
                           a(3) => N309, a(2) => N308, a(1) => N307, a(0) => 
                           n18, b(31) => net35534, b(30) => net35534, b(29) => 
                           net35534, b(28) => net35534, b(27) => net35534, 
                           b(26) => net35534, b(25) => net35534, b(24) => 
                           net35534, b(23) => net35534, b(22) => net35534, 
                           b(21) => net35534, b(20) => net35534, b(19) => 
                           net35534, b(18) => net35534, b(17) => net35534, 
                           b(16) => net35534, b(15) => net35534, b(14) => 
                           net35534, b(13) => net35534, b(12) => net35534, 
                           b(11) => net35534, b(10) => net35534, b(9) => 
                           net35534, b(8) => net35534, b(7) => net35534, b(6) 
                           => net35534, b(5) => net35534, b(4) => net35534, 
                           b(3) => net35534, b(2) => n7, b(1) => n7, b(0) => n7
                           , quotient(4) => n_1724, quotient(3) => n_1725, 
                           quotient(2) => n_1726, quotient(1) => n_1727, 
                           quotient(0) => n_1728, remainder(31) => n_1729, 
                           remainder(30) => n_1730, remainder(29) => n_1731, 
                           remainder(28) => n_1732, remainder(27) => n_1733, 
                           remainder(26) => n_1734, remainder(25) => n_1735, 
                           remainder(24) => n_1736, remainder(23) => n_1737, 
                           remainder(22) => n_1738, remainder(21) => n_1739, 
                           remainder(20) => n_1740, remainder(19) => n_1741, 
                           remainder(18) => n_1742, remainder(17) => n_1743, 
                           remainder(16) => n_1744, remainder(15) => n_1745, 
                           remainder(14) => n_1746, remainder(13) => n_1747, 
                           remainder(12) => n_1748, remainder(11) => n_1749, 
                           remainder(10) => n_1750, remainder(9) => n_1751, 
                           remainder(8) => n_1752, remainder(7) => n_1753, 
                           remainder(6) => n_1754, remainder(5) => n_1755, 
                           remainder(4) => n_1756, remainder(3) => n_1757, 
                           remainder(2) => N2, remainder(1) => N1, remainder(0)
                           => N0, divide_by_0 => n_1723);
   add_219_2_U1_1_1 : HAxp5_ASAP7_75t_R port map( A => crossbar_ctrl_vec(1), B 
                           => crossbar_ctrl_vec(0), CON => n23, SN => n22);
   add_219_2_U1_1_2 : HAxp5_ASAP7_75t_R port map( A => crossbar_ctrl_vec(2), B 
                           => n26, CON => n25, SN => n24);
   U3 : XOR2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_8_port, B => n4, Y => 
                           n1_port);
   U4 : XNOR2xp5_ASAP7_75t_R port map( A => n8, B => crossbar_ctrl_14_port, Y 
                           => n2_port);
   U5 : XNOR2xp5_ASAP7_75t_R port map( A => n6, B => crossbar_ctrl_20_port, Y 
                           => n3);
   U6 : OR2x2_ASAP7_75t_R port map( A => crossbar_ctrl_6_port, B => 
                           crossbar_ctrl_7_port, Y => n4);
   U7 : XOR2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_5_port, B => 
                           crossbar_ctrl_4_port, Y => n5);
   U8 : OR2x2_ASAP7_75t_R port map( A => crossbar_ctrl_18_port, B => 
                           crossbar_ctrl_19_port, Y => n6);
   U9 : AND2x2_ASAP7_75t_R port map( A => crossbar_ctrl_13_port, B => 
                           crossbar_ctrl_12_port, Y => n8);
   U10 : XNOR2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_6_port, B => 
                           crossbar_ctrl_7_port, Y => n9);
   U11 : AND2x2_ASAP7_75t_R port map( A => crossbar_ctrl_8_port, B => n4, Y => 
                           n10);
   U12 : XNOR2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_16_port, B => 
                           crossbar_ctrl_17_port, Y => n11);
   U13 : AND2x2_ASAP7_75t_R port map( A => crossbar_ctrl_5_port, B => 
                           crossbar_ctrl_4_port, Y => n12);
   U14 : OR2x2_ASAP7_75t_R port map( A => n6, B => crossbar_ctrl_20_port, Y => 
                           n13);
   U15 : XNOR2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_18_port, B => 
                           crossbar_ctrl_19_port, Y => n14);
   U16 : XOR2xp5_ASAP7_75t_R port map( A => crossbar_ctrl_13_port, B => 
                           crossbar_ctrl_12_port, Y => n15);
   U17 : OR2x2_ASAP7_75t_R port map( A => crossbar_ctrl_16_port, B => 
                           crossbar_ctrl_17_port, Y => n16);
   U18 : OR2x2_ASAP7_75t_R port map( A => n8, B => crossbar_ctrl_14_port, Y => 
                           n17);
   U19 : NOR2xp33_ASAP7_75t_R port map( A => n29, B => n72, Y => 
                           vc_transfer_vec(10));
   U20 : NOR2xp33_ASAP7_75t_R port map( A => n52, B => n127, Y => n113);
   U21 : NOR2xp33_ASAP7_75t_R port map( A => n29, B => n73, Y => 
                           vc_transfer_vec(9));
   U22 : NOR2xp33_ASAP7_75t_R port map( A => n37, B => n122, Y => n109);
   U23 : NOR2xp33_ASAP7_75t_R port map( A => n40, B => n121, Y => n110);
   U24 : NOR2xp33_ASAP7_75t_R port map( A => n43, B => n123, Y => n108);
   U25 : NOR2xp33_ASAP7_75t_R port map( A => n49, B => n124, Y => n112);
   U26 : NOR2xp33_ASAP7_75t_R port map( A => n28, B => n69, Y => 
                           vc_transfer_vec(8));
   U27 : NOR2xp33_ASAP7_75t_R port map( A => n28, B => n70, Y => 
                           vc_transfer_vec(7));
   U28 : NOR2xp33_ASAP7_75t_R port map( A => n33_port, B => n61, Y => 
                           vc_transfer_vec(4));
   U29 : NOR2xp33_ASAP7_75t_R port map( A => n33_port, B => n63, Y => 
                           vc_transfer_vec(3));
   U30 : NOR2xp33_ASAP7_75t_R port map( A => n127, B => N194, Y => n103);
   U31 : NOR2xp33_ASAP7_75t_R port map( A => n122, B => N34, Y => n99);
   U32 : NOR2xp33_ASAP7_75t_R port map( A => n46, B => n125, Y => n111);
   U33 : NOR2xp33_ASAP7_75t_R port map( A => n123, B => N98, Y => n98_port);
   U34 : NOR2xp33_ASAP7_75t_R port map( A => n121, B => N66, Y => n100);
   U36 : NOR2xp33_ASAP7_75t_R port map( A => n124, B => N162, Y => n102);
   U39 : NOR2xp33_ASAP7_75t_R port map( A => n31, B => n74, Y => 
                           vc_transfer_vec(12));
   U44 : NOR2xp33_ASAP7_75t_R port map( A => n125, B => N130, Y => n101);
   U45 : NOR2xp33_ASAP7_75t_R port map( A => n27, B => n56, Y => 
                           vc_transfer_vec(2));
   U46 : NOR2xp33_ASAP7_75t_R port map( A => n32_port, B => n66_port, Y => 
                           vc_transfer_vec(6));
   U47 : NOR2xp33_ASAP7_75t_R port map( A => n32_port, B => n67, Y => 
                           vc_transfer_vec(5));
   U50 : NOR2xp33_ASAP7_75t_R port map( A => n31, B => n75, Y => 
                           vc_transfer_vec(11));
   U53 : NOR2xp33_ASAP7_75t_R port map( A => n27, B => n59, Y => 
                           vc_transfer_vec(1));
   U54 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec(0), B => 
                           n66_port, Y => n150);
   U61 : NOR2xp33_ASAP7_75t_R port map( A => n72, B => n248, Y => n221);
   U62 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_18_port, Y => n19);
   U63 : NOR2xp33_ASAP7_75t_R port map( A => n72, B => n246, Y => n225);
   U66 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(0), Y => n18);
   U67 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx_vec_5_port, B => 
                           vc_write_tx_vec_6_port, Y => n123);
   U68 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx_vec_1_port, B => 
                           vc_write_tx_vec_2_port, Y => n122);
   U79 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx_vec_10_port, B => 
                           vc_write_tx_vec_9_port, Y => n124);
   U80 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx_vec_3_port, B => 
                           vc_write_tx_vec_4_port, Y => n121);
   U81 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx_vec_11_port, B => 
                           vc_write_tx_vec_12_port, Y => n127);
   U84 : NOR2xp33_ASAP7_75t_R port map( A => vc_write_tx_vec_7_port, B => 
                           vc_write_tx_vec_8_port, Y => n125);
   U85 : AOI31xp33_ASAP7_75t_R port map( A1 => n94, A2 => n95, A3 => n96_port, 
                           B => n97_port, Y => vc_transfer_vec(0));
   U86 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec(30), B => n67, Y
                           => n235);
   U87 : INVx1_ASAP7_75t_R port map( A => n97_port, Y => n249);
   U90 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec(18), B => n56, Y
                           => n181);
   U91 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec(27), B => n75, Y
                           => n160_port);
   U94 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec(15), B => n56, Y
                           => n191);
   U97 : NOR2xp33_ASAP7_75t_R port map( A => n126, B => N2, Y => n104);
   U100 : NOR2xp33_ASAP7_75t_R port map( A => n245, B => n220, Y => 
                           channel_rq_12_port);
   U101 : NOR3xp33_ASAP7_75t_R port map( A => n253, B => crossbar_ctrl_vec(8), 
                           C => n67, Y => n205);
   U114 : NOR3xp33_ASAP7_75t_R port map( A => n84, B => crossbar_ctrl_vec(19), 
                           C => n73, Y => n177);
   U115 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec(6), B => n69, Y
                           => n209);
   U116 : NOR3xp33_ASAP7_75t_R port map( A => n84, B => crossbar_ctrl_vec(19), 
                           C => n72, Y => n180);
   U117 : NOR2xp33_ASAP7_75t_R port map( A => n247, B => n224, Y => 
                           channel_rq_11_port);
   U118 : NOR3xp33_ASAP7_75t_R port map( A => n250, B => crossbar_ctrl_vec(5), 
                           C => n67, Y => n215);
   U119 : NOR3xp33_ASAP7_75t_R port map( A => n253, B => crossbar_ctrl_vec(8), 
                           C => n66_port, Y => n208);
   U120 : NOR3xp33_ASAP7_75t_R port map( A => n81, B => crossbar_ctrl_vec(16), 
                           C => n73, Y => n187);
   U121 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec(32), B => 
                           crossbar_ctrl_vec(31), Y => n237);
   U122 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec(30), B => n75, 
                           Y => n236);
   U123 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec(3), B => n69, Y
                           => n219);
   U124 : NOR3xp33_ASAP7_75t_R port map( A => n81, B => crossbar_ctrl_vec(16), 
                           C => n72, Y => n190);
   U125 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec(27), B => n67, 
                           Y => n159);
   U126 : NOR3xp33_ASAP7_75t_R port map( A => n250, B => crossbar_ctrl_vec(5), 
                           C => n66_port, Y => n218);
   U127 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec(29), B => 
                           crossbar_ctrl_vec(28), Y => n161_port);
   U128 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec(0), B => n72, Y
                           => n151);
   U129 : NOR2xp33_ASAP7_75t_R port map( A => crossbar_ctrl_vec(0), B => n56, Y
                           => n145);
   U130 : NOR3xp33_ASAP7_75t_R port map( A => n144, B => crossbar_ctrl_vec(2), 
                           C => crossbar_ctrl_vec(1), Y => n143);
   U131 : HB1xp67_ASAP7_75t_R port map( A => rst, Y => n20);
   U132 : HB1xp67_ASAP7_75t_R port map( A => rst, Y => n21);
   U133 : TIEHIx1_ASAP7_75t_R port map( H => n7);
   U134 : TIELOx1_ASAP7_75t_R port map( L => net35534);
   U135 : INVx1_ASAP7_75t_R port map( A => n22, Y => N307);
   U136 : INVx1_ASAP7_75t_R port map( A => n23, Y => n26);
   U137 : INVx1_ASAP7_75t_R port map( A => n24, Y => N308);
   U138 : INVx1_ASAP7_75t_R port map( A => n25, Y => N309);
   U139 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_4_port, Y => N330);
   U140 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_6_port, Y => N353);
   U141 : INVx1_ASAP7_75t_R port map( A => N380, Y => N379);
   U142 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_12_port, Y => N401);
   U143 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_16_port, Y => N426);
   U144 : INVx1_ASAP7_75t_R port map( A => switch_ack_var_1_port, Y => n27);
   U145 : INVx1_ASAP7_75t_R port map( A => switch_ack_var_4_port, Y => n28);
   U146 : INVx1_ASAP7_75t_R port map( A => switch_ack_var_5_port, Y => n29);
   U147 : INVx1_ASAP7_75t_R port map( A => N1, Y => n30);
   U148 : INVx1_ASAP7_75t_R port map( A => switch_ack_var_6_port, Y => n31);
   U149 : INVx1_ASAP7_75t_R port map( A => switch_ack_var_3_port, Y => n32_port
                           );
   U150 : INVx1_ASAP7_75t_R port map( A => switch_ack_var_2_port, Y => n33_port
                           );
   U151 : INVx1_ASAP7_75t_R port map( A => N0, Y => n34_port);
   U152 : INVx1_ASAP7_75t_R port map( A => N33, Y => n35);
   U153 : INVx1_ASAP7_75t_R port map( A => N32, Y => n36);
   U154 : INVx1_ASAP7_75t_R port map( A => N34, Y => n37);
   U155 : INVx1_ASAP7_75t_R port map( A => N65, Y => n38);
   U156 : INVx1_ASAP7_75t_R port map( A => N64, Y => n39);
   U157 : INVx1_ASAP7_75t_R port map( A => N66, Y => n40);
   U158 : INVx1_ASAP7_75t_R port map( A => N97, Y => n41);
   U159 : INVx1_ASAP7_75t_R port map( A => N96, Y => n42);
   U160 : INVx1_ASAP7_75t_R port map( A => N98, Y => n43);
   U161 : INVx1_ASAP7_75t_R port map( A => N129, Y => n44);
   U162 : INVx1_ASAP7_75t_R port map( A => N128, Y => n45);
   U163 : INVx1_ASAP7_75t_R port map( A => N130, Y => n46);
   U164 : INVx1_ASAP7_75t_R port map( A => N161, Y => n47);
   U165 : INVx1_ASAP7_75t_R port map( A => N160, Y => n48);
   U166 : INVx1_ASAP7_75t_R port map( A => N162, Y => n49);
   U167 : INVx1_ASAP7_75t_R port map( A => N193, Y => n50);
   U168 : INVx1_ASAP7_75t_R port map( A => N192, Y => n51);
   U169 : INVx1_ASAP7_75t_R port map( A => N194, Y => n52);
   U170 : INVx1_ASAP7_75t_R port map( A => vc_write_tx_vec_9_port, Y => n53);
   U171 : INVx1_ASAP7_75t_R port map( A => n126, Y => vc_write_tx_vec_0_port);
   U172 : INVx1_ASAP7_75t_R port map( A => vc_write_tx_vec_5_port, Y => n55);
   U173 : INVx1_ASAP7_75t_R port map( A => poss_channel_rq_5_2_1_port, Y => n56
                           );
   U174 : INVx1_ASAP7_75t_R port map( A => n176, Y => n57);
   U175 : INVx1_ASAP7_75t_R port map( A => n186, Y => n58);
   U176 : INVx1_ASAP7_75t_R port map( A => poss_channel_rq_5_2_0_port, Y => n59
                           );
   U177 : INVx1_ASAP7_75t_R port map( A => vc_write_tx_vec_7_port, Y => n60);
   U178 : INVx1_ASAP7_75t_R port map( A => poss_channel_rq_5_3_1_port, Y => n61
                           );
   U179 : INVx1_ASAP7_75t_R port map( A => vc_write_tx_vec_1_port, Y => n62);
   U180 : INVx1_ASAP7_75t_R port map( A => poss_channel_rq_5_3_0_port, Y => n63
                           );
   U181 : INVx1_ASAP7_75t_R port map( A => n204, Y => n64_port);
   U182 : INVx1_ASAP7_75t_R port map( A => n214, Y => n65_port);
   U183 : INVx1_ASAP7_75t_R port map( A => poss_channel_rq_5_4_1_port, Y => 
                           n66_port);
   U184 : INVx1_ASAP7_75t_R port map( A => poss_channel_rq_5_4_0_port, Y => n67
                           );
   U185 : INVx1_ASAP7_75t_R port map( A => vc_write_tx_vec_3_port, Y => n68);
   U186 : INVx1_ASAP7_75t_R port map( A => poss_channel_rq_5_5_1_port, Y => n69
                           );
   U187 : INVx1_ASAP7_75t_R port map( A => poss_channel_rq_5_5_0_port, Y => n70
                           );
   U188 : INVx1_ASAP7_75t_R port map( A => vc_write_tx_vec_11_port, Y => n71);
   U189 : INVx1_ASAP7_75t_R port map( A => poss_channel_rq_6_5_1_port, Y => n72
                           );
   U190 : INVx1_ASAP7_75t_R port map( A => poss_channel_rq_6_5_0_port, Y => n73
                           );
   U191 : INVx1_ASAP7_75t_R port map( A => poss_channel_rq_5_0_1_port, Y => n74
                           );
   U192 : INVx1_ASAP7_75t_R port map( A => poss_channel_rq_5_0_0_port, Y => n75
                           );
   U193 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(9), Y => n76);
   U194 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_vec(3), Y => n77);
   U195 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(12), Y => n78);
   U196 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(13), Y => n79);
   U197 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_vec(4), Y => n80);
   U198 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(15), Y => n81);
   U199 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(17), Y => n82);
   U298 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_vec(5), Y => n83);
   U299 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(18), Y => n84);
   U300 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(20), Y => n85);
   U301 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_vec(6), Y => n86);
   U302 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(22), Y => n87);
   U303 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(23), Y => n88);
   U304 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_vec(7), Y => n89);
   U305 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(25), Y => n90);
   U306 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(26), Y => n91);
   U307 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_vec(8), Y => n92);
   U308 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(27), Y => n93);
   U309 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(28), Y => n240);
   U310 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(29), Y => n241);
   U311 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(30), Y => n242);
   U312 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(31), Y => n243);
   U313 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(32), Y => n244);
   U314 : INVx1_ASAP7_75t_R port map( A => output_vc_in_use(12), Y => n245);
   U315 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(33), Y => n246);
   U316 : INVx1_ASAP7_75t_R port map( A => output_vc_in_use(11), Y => n247);
   U317 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(36), Y => n248);
   U318 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(3), Y => n250);
   U319 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(4), Y => n251);
   U320 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_vec(1), Y => n252);
   U321 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(6), Y => n253);
   U322 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(7), Y => n254);
   U323 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_vec(2), Y => n255);
   U324 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(2), Y => n256);
   U325 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl_vec(1), Y => n257);
   U326 : INVx1_ASAP7_75t_R port map( A => vc_sel_enc_vec(0), Y => n258);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity vc_allocator_7_1_1_1_1_DXYU is

   port( clk, rst : in std_logic;  header : in std_logic_vector (129 downto 0);
         enr_vc, valid_data_vc_vec : in std_logic_vector (12 downto 0);  
         input_vc_in_use : out std_logic_vector (12 downto 0);  
         crossbar_ctrl_vec : out std_logic_vector (38 downto 0);  
         vc_sel_enc_vec, output_vc_in_use : out std_logic_vector (12 downto 0)
         );

end vc_allocator_7_1_1_1_1_DXYU;

architecture SYN_rtl of vc_allocator_7_1_1_1_1_DXYU is

   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component vc_output_allocator_port_num7_vc_num_out2_1
      port( clk, rst : in std_logic;  rq_vc_out : in std_logic_vector (5 downto
            0);  granted_vc, packet_end : in std_logic_vector (11 downto 0);  
            crossbar_ctrl_vec : out std_logic_vector (5 downto 0);  vc_sel_enc,
            output_vc_in_use : out std_logic_vector (1 downto 0);  
            ack_rq_vc_out : out std_logic_vector (5 downto 0));
   end component;
   
   component header_arbiter_and_decoder_1_1_1_7_6_2_1_DXYU
      port( clk, rst : in std_logic;  header : in std_logic_vector (19 downto 
            0);  valid_data_vc, enr_vc : in std_logic_vector (1 downto 0);  
            ack_vc : in std_logic;  granted_rq : out std_logic_vector (6 downto
            0);  input_vc_in_use, packet_end, granted_vc : out std_logic_vector
            (1 downto 0));
   end component;
   
   component vc_output_allocator_port_num7_vc_num_out2_2
      port( clk, rst : in std_logic;  rq_vc_out : in std_logic_vector (5 downto
            0);  granted_vc, packet_end : in std_logic_vector (11 downto 0);  
            crossbar_ctrl_vec : out std_logic_vector (5 downto 0);  vc_sel_enc,
            output_vc_in_use : out std_logic_vector (1 downto 0);  
            ack_rq_vc_out : out std_logic_vector (5 downto 0));
   end component;
   
   component header_arbiter_and_decoder_1_1_1_7_5_2_1_DXYU
      port( clk, rst : in std_logic;  header : in std_logic_vector (19 downto 
            0);  valid_data_vc, enr_vc : in std_logic_vector (1 downto 0);  
            ack_vc : in std_logic;  granted_rq : out std_logic_vector (6 downto
            0);  input_vc_in_use, packet_end, granted_vc : out std_logic_vector
            (1 downto 0));
   end component;
   
   component vc_output_allocator_port_num7_vc_num_out2_3
      port( clk, rst : in std_logic;  rq_vc_out : in std_logic_vector (5 downto
            0);  granted_vc, packet_end : in std_logic_vector (11 downto 0);  
            crossbar_ctrl_vec : out std_logic_vector (5 downto 0);  vc_sel_enc,
            output_vc_in_use : out std_logic_vector (1 downto 0);  
            ack_rq_vc_out : out std_logic_vector (5 downto 0));
   end component;
   
   component header_arbiter_and_decoder_1_1_1_7_4_2_1_DXYU
      port( clk, rst : in std_logic;  header : in std_logic_vector (19 downto 
            0);  valid_data_vc, enr_vc : in std_logic_vector (1 downto 0);  
            ack_vc : in std_logic;  granted_rq : out std_logic_vector (6 downto
            0);  input_vc_in_use, packet_end, granted_vc : out std_logic_vector
            (1 downto 0));
   end component;
   
   component vc_output_allocator_port_num7_vc_num_out2_4
      port( clk, rst : in std_logic;  rq_vc_out : in std_logic_vector (5 downto
            0);  granted_vc, packet_end : in std_logic_vector (11 downto 0);  
            crossbar_ctrl_vec : out std_logic_vector (5 downto 0);  vc_sel_enc,
            output_vc_in_use : out std_logic_vector (1 downto 0);  
            ack_rq_vc_out : out std_logic_vector (5 downto 0));
   end component;
   
   component header_arbiter_and_decoder_1_1_1_7_3_2_1_DXYU
      port( clk, rst : in std_logic;  header : in std_logic_vector (19 downto 
            0);  valid_data_vc, enr_vc : in std_logic_vector (1 downto 0);  
            ack_vc : in std_logic;  granted_rq : out std_logic_vector (6 downto
            0);  input_vc_in_use, packet_end, granted_vc : out std_logic_vector
            (1 downto 0));
   end component;
   
   component vc_output_allocator_port_num7_vc_num_out2_5
      port( clk, rst : in std_logic;  rq_vc_out : in std_logic_vector (5 downto
            0);  granted_vc, packet_end : in std_logic_vector (11 downto 0);  
            crossbar_ctrl_vec : out std_logic_vector (5 downto 0);  vc_sel_enc,
            output_vc_in_use : out std_logic_vector (1 downto 0);  
            ack_rq_vc_out : out std_logic_vector (5 downto 0));
   end component;
   
   component header_arbiter_and_decoder_1_1_1_7_2_2_1_DXYU
      port( clk, rst : in std_logic;  header : in std_logic_vector (19 downto 
            0);  valid_data_vc, enr_vc : in std_logic_vector (1 downto 0);  
            ack_vc : in std_logic;  granted_rq : out std_logic_vector (6 downto
            0);  input_vc_in_use, packet_end, granted_vc : out std_logic_vector
            (1 downto 0));
   end component;
   
   component vc_output_allocator_port_num7_vc_num_out2_0
      port( clk, rst : in std_logic;  rq_vc_out : in std_logic_vector (5 downto
            0);  granted_vc, packet_end : in std_logic_vector (11 downto 0);  
            crossbar_ctrl_vec : out std_logic_vector (5 downto 0);  vc_sel_enc,
            output_vc_in_use : out std_logic_vector (1 downto 0);  
            ack_rq_vc_out : out std_logic_vector (5 downto 0));
   end component;
   
   component header_arbiter_and_decoder_1_1_1_7_1_2_1_DXYU
      port( clk, rst : in std_logic;  header : in std_logic_vector (19 downto 
            0);  valid_data_vc, enr_vc : in std_logic_vector (1 downto 0);  
            ack_vc : in std_logic;  granted_rq : out std_logic_vector (6 downto
            0);  input_vc_in_use, packet_end, granted_vc : out std_logic_vector
            (1 downto 0));
   end component;
   
   component vc_output_allocator_port_num7_vc_num_out1
      port( clk, rst : in std_logic;  rq_vc_out : in std_logic_vector (5 downto
            0);  granted_vc, packet_end : in std_logic_vector (11 downto 0);  
            crossbar_ctrl_vec : out std_logic_vector (2 downto 0);  vc_sel_enc,
            output_vc_in_use : out std_logic;  ack_rq_vc_out : out 
            std_logic_vector (5 downto 0));
   end component;
   
   component header_arbiter_and_decoder_1_1_1_7_0_1_1_DXYU
      port( clk, rst : in std_logic;  header : in std_logic_vector (9 downto 0)
            ;  valid_data_vc, enr_vc, ack_vc : in std_logic;  granted_rq : out 
            std_logic_vector (6 downto 0);  input_vc_in_use, packet_end, 
            granted_vc : out std_logic);
   end component;
   
   component OR3x1_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR4x1_ASAP7_75t_R
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OR5x1_ASAP7_75t_R
      port( A, B, C, D, E : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2x2_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic0_port, ack_rq_vc_out_6_5_port, ack_rq_vc_out_6_0_port, 
      ack_rq_vc_out_5_5_port, ack_rq_vc_out_5_4_port, ack_rq_vc_out_5_3_port, 
      ack_rq_vc_out_5_2_port, ack_rq_vc_out_5_1_port, ack_rq_vc_out_5_0_port, 
      ack_rq_vc_out_4_4_port, ack_rq_vc_out_4_2_port, ack_rq_vc_out_4_0_port, 
      ack_rq_vc_out_3_5_port, ack_rq_vc_out_3_4_port, ack_rq_vc_out_3_3_port, 
      ack_rq_vc_out_3_1_port, ack_rq_vc_out_3_0_port, ack_rq_vc_out_2_4_port, 
      ack_rq_vc_out_2_2_port, ack_rq_vc_out_2_1_port, ack_rq_vc_out_1_5_port, 
      ack_rq_vc_out_1_3_port, ack_rq_vc_out_1_2_port, ack_rq_vc_out_1_1_port, 
      ack_rq_vc_out_1_0_port, ack_rq_vc_out_0_5_port, ack_rq_vc_out_0_4_port, 
      ack_rq_vc_out_0_3_port, ack_rq_vc_out_0_2_port, ack_rq_vc_out_0_1_port, 
      ack_rq_vc_out_0_0_port, packet_end_sort_6_5_1_port, 
      packet_end_sort_6_5_0_port, packet_end_sort_6_0_0_port, 
      packet_end_sort_5_5_1_port, packet_end_sort_5_5_0_port, 
      packet_end_sort_5_4_1_port, packet_end_sort_5_4_0_port, 
      packet_end_sort_5_3_1_port, packet_end_sort_5_3_0_port, 
      packet_end_sort_5_2_1_port, packet_end_sort_5_2_0_port, 
      packet_end_sort_5_0_1_port, packet_end_sort_5_0_0_port, 
      granted_vc_sort_6_5_1_port, granted_vc_sort_6_5_0_port, 
      granted_vc_sort_6_0_0_port, granted_vc_sort_5_5_1_port, 
      granted_vc_sort_5_5_0_port, granted_vc_sort_5_4_1_port, 
      granted_vc_sort_5_4_0_port, granted_vc_sort_5_3_1_port, 
      granted_vc_sort_5_3_0_port, granted_vc_sort_5_2_1_port, 
      granted_vc_sort_5_2_0_port, granted_vc_sort_5_0_1_port, 
      granted_vc_sort_5_0_0_port, rq_vc_out_array_6_5_port, 
      rq_vc_out_array_6_0_port, rq_vc_out_array_5_5_port, 
      rq_vc_out_array_5_4_port, rq_vc_out_array_5_3_port, 
      rq_vc_out_array_5_2_port, rq_vc_out_array_5_1_port, 
      rq_vc_out_array_5_0_port, rq_vc_out_array_4_4_port, 
      rq_vc_out_array_4_2_port, rq_vc_out_array_4_0_port, 
      rq_vc_out_array_3_5_port, rq_vc_out_array_3_4_port, 
      rq_vc_out_array_3_3_port, rq_vc_out_array_3_1_port, 
      rq_vc_out_array_3_0_port, rq_vc_out_array_2_4_port, 
      rq_vc_out_array_2_2_port, rq_vc_out_array_2_1_port, 
      rq_vc_out_array_1_5_port, rq_vc_out_array_1_3_port, 
      rq_vc_out_array_1_2_port, rq_vc_out_array_1_1_port, 
      rq_vc_out_array_1_0_port, rq_vc_out_array_0_5_port, 
      rq_vc_out_array_0_4_port, rq_vc_out_array_0_3_port, 
      rq_vc_out_array_0_2_port, rq_vc_out_array_0_1_port, 
      rq_vc_out_array_0_0_port, ack_rq_vc_out_var_6_port, 
      ack_rq_vc_out_var_5_port, ack_rq_vc_out_var_4_port, 
      ack_rq_vc_out_var_3_port, ack_rq_vc_out_var_2_port, 
      ack_rq_vc_out_var_1_port, ack_rq_vc_out_var_0_port, n1, n2, n3, n_1758, 
      n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, 
      n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, 
      n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, 
      n_1786, n_1787, n_1788 : std_logic;

begin
   
   U2 : OR2x2_ASAP7_75t_R port map( A => ack_rq_vc_out_0_5_port, B => 
                           ack_rq_vc_out_5_0_port, Y => 
                           ack_rq_vc_out_var_6_port);
   U3 : OR4x1_ASAP7_75t_R port map( A => ack_rq_vc_out_2_2_port, B => 
                           ack_rq_vc_out_1_3_port, C => ack_rq_vc_out_0_4_port,
                           D => n1, Y => ack_rq_vc_out_var_5_port);
   U4 : OR3x1_ASAP7_75t_R port map( A => ack_rq_vc_out_6_5_port, B => 
                           ack_rq_vc_out_4_0_port, C => ack_rq_vc_out_3_1_port,
                           Y => n1);
   U5 : OR5x1_ASAP7_75t_R port map( A => ack_rq_vc_out_5_5_port, B => 
                           ack_rq_vc_out_3_0_port, C => ack_rq_vc_out_2_1_port,
                           D => ack_rq_vc_out_1_2_port, E => 
                           ack_rq_vc_out_0_3_port, Y => 
                           ack_rq_vc_out_var_4_port);
   U6 : OR3x1_ASAP7_75t_R port map( A => ack_rq_vc_out_5_4_port, B => 
                           ack_rq_vc_out_1_1_port, C => ack_rq_vc_out_0_2_port,
                           Y => ack_rq_vc_out_var_3_port);
   U7 : OR5x1_ASAP7_75t_R port map( A => ack_rq_vc_out_5_3_port, B => 
                           ack_rq_vc_out_4_4_port, C => ack_rq_vc_out_3_5_port,
                           D => ack_rq_vc_out_1_0_port, E => 
                           ack_rq_vc_out_0_1_port, Y => 
                           ack_rq_vc_out_var_2_port);
   U8 : OR3x1_ASAP7_75t_R port map( A => ack_rq_vc_out_5_2_port, B => 
                           ack_rq_vc_out_3_4_port, C => ack_rq_vc_out_0_0_port,
                           Y => ack_rq_vc_out_var_1_port);
   U9 : OR4x1_ASAP7_75t_R port map( A => ack_rq_vc_out_3_3_port, B => 
                           ack_rq_vc_out_2_4_port, C => ack_rq_vc_out_1_5_port,
                           D => n2, Y => ack_rq_vc_out_var_0_port);
   U10 : OR3x1_ASAP7_75t_R port map( A => ack_rq_vc_out_6_0_port, B => 
                           ack_rq_vc_out_5_1_port, C => ack_rq_vc_out_4_2_port,
                           Y => n2);
   input_first_arbiter_i_0 : header_arbiter_and_decoder_1_1_1_7_0_1_1_DXYU port
                           map( clk => clk, rst => n3, header(9) => header(9), 
                           header(8) => header(8), header(7) => header(7), 
                           header(6) => header(6), header(5) => header(5), 
                           header(4) => header(4), header(3) => header(3), 
                           header(2) => header(2), header(1) => header(1), 
                           header(0) => header(0), valid_data_vc => 
                           valid_data_vc_vec(0), enr_vc => enr_vc(0), ack_vc =>
                           ack_rq_vc_out_var_0_port, granted_rq(6) => 
                           rq_vc_out_array_6_0_port, granted_rq(5) => 
                           rq_vc_out_array_5_1_port, granted_rq(4) => 
                           rq_vc_out_array_4_2_port, granted_rq(3) => 
                           rq_vc_out_array_3_3_port, granted_rq(2) => 
                           rq_vc_out_array_2_4_port, granted_rq(1) => 
                           rq_vc_out_array_1_5_port, granted_rq(0) => n_1758, 
                           input_vc_in_use => input_vc_in_use(0), packet_end =>
                           packet_end_sort_6_0_0_port, granted_vc => 
                           granted_vc_sort_6_0_0_port);
   output_last_arbiter_i_0 : vc_output_allocator_port_num7_vc_num_out1 port 
                           map( clk => clk, rst => n3, rq_vc_out(5) => 
                           rq_vc_out_array_0_5_port, rq_vc_out(4) => 
                           rq_vc_out_array_0_4_port, rq_vc_out(3) => 
                           rq_vc_out_array_0_3_port, rq_vc_out(2) => 
                           rq_vc_out_array_0_2_port, rq_vc_out(1) => 
                           rq_vc_out_array_0_1_port, rq_vc_out(0) => 
                           rq_vc_out_array_0_0_port, granted_vc(11) => 
                           granted_vc_sort_5_0_1_port, granted_vc(10) => 
                           granted_vc_sort_5_0_0_port, granted_vc(9) => 
                           granted_vc_sort_6_5_1_port, granted_vc(8) => 
                           granted_vc_sort_6_5_0_port, granted_vc(7) => 
                           granted_vc_sort_5_5_1_port, granted_vc(6) => 
                           granted_vc_sort_5_5_0_port, granted_vc(5) => 
                           granted_vc_sort_5_4_1_port, granted_vc(4) => 
                           granted_vc_sort_5_4_0_port, granted_vc(3) => 
                           granted_vc_sort_5_3_1_port, granted_vc(2) => 
                           granted_vc_sort_5_3_0_port, granted_vc(1) => 
                           granted_vc_sort_5_2_1_port, granted_vc(0) => 
                           granted_vc_sort_5_2_0_port, packet_end(11) => 
                           packet_end_sort_5_0_1_port, packet_end(10) => 
                           packet_end_sort_5_0_0_port, packet_end(9) => 
                           packet_end_sort_6_5_1_port, packet_end(8) => 
                           packet_end_sort_6_5_0_port, packet_end(7) => 
                           packet_end_sort_5_5_1_port, packet_end(6) => 
                           packet_end_sort_5_5_0_port, packet_end(5) => 
                           packet_end_sort_5_4_1_port, packet_end(4) => 
                           packet_end_sort_5_4_0_port, packet_end(3) => 
                           packet_end_sort_5_3_1_port, packet_end(2) => 
                           packet_end_sort_5_3_0_port, packet_end(1) => 
                           packet_end_sort_5_2_1_port, packet_end(0) => 
                           packet_end_sort_5_2_0_port, crossbar_ctrl_vec(2) => 
                           crossbar_ctrl_vec(2), crossbar_ctrl_vec(1) => 
                           crossbar_ctrl_vec(1), crossbar_ctrl_vec(0) => 
                           crossbar_ctrl_vec(0), vc_sel_enc => 
                           vc_sel_enc_vec(0), output_vc_in_use => 
                           output_vc_in_use(0), ack_rq_vc_out(5) => 
                           ack_rq_vc_out_0_5_port, ack_rq_vc_out(4) => 
                           ack_rq_vc_out_0_4_port, ack_rq_vc_out(3) => 
                           ack_rq_vc_out_0_3_port, ack_rq_vc_out(2) => 
                           ack_rq_vc_out_0_2_port, ack_rq_vc_out(1) => 
                           ack_rq_vc_out_0_1_port, ack_rq_vc_out(0) => 
                           ack_rq_vc_out_0_0_port);
   input_first_arbiter_i_1 : header_arbiter_and_decoder_1_1_1_7_1_2_1_DXYU port
                           map( clk => clk, rst => n3, header(19) => header(29)
                           , header(18) => header(28), header(17) => header(27)
                           , header(16) => header(26), header(15) => header(25)
                           , header(14) => header(24), header(13) => header(23)
                           , header(12) => header(22), header(11) => header(21)
                           , header(10) => header(20), header(9) => header(19),
                           header(8) => header(18), header(7) => header(17), 
                           header(6) => header(16), header(5) => header(15), 
                           header(4) => header(14), header(3) => header(13), 
                           header(2) => header(12), header(1) => header(11), 
                           header(0) => header(10), valid_data_vc(1) => 
                           valid_data_vc_vec(2), valid_data_vc(0) => 
                           valid_data_vc_vec(1), enr_vc(1) => enr_vc(2), 
                           enr_vc(0) => enr_vc(1), ack_vc => 
                           ack_rq_vc_out_var_1_port, granted_rq(6) => n_1759, 
                           granted_rq(5) => rq_vc_out_array_5_2_port, 
                           granted_rq(4) => n_1760, granted_rq(3) => 
                           rq_vc_out_array_3_4_port, granted_rq(2) => n_1761, 
                           granted_rq(1) => n_1762, granted_rq(0) => 
                           rq_vc_out_array_0_0_port, input_vc_in_use(1) => 
                           input_vc_in_use(2), input_vc_in_use(0) => 
                           input_vc_in_use(1), packet_end(1) => 
                           packet_end_sort_5_2_1_port, packet_end(0) => 
                           packet_end_sort_5_2_0_port, granted_vc(1) => 
                           granted_vc_sort_5_2_1_port, granted_vc(0) => 
                           granted_vc_sort_5_2_0_port);
   output_last_arbiter_i_1 : vc_output_allocator_port_num7_vc_num_out2_0 port 
                           map( clk => clk, rst => n3, rq_vc_out(5) => 
                           rq_vc_out_array_1_5_port, rq_vc_out(4) => 
                           X_Logic0_port, rq_vc_out(3) => 
                           rq_vc_out_array_1_3_port, rq_vc_out(2) => 
                           rq_vc_out_array_1_2_port, rq_vc_out(1) => 
                           rq_vc_out_array_1_1_port, rq_vc_out(0) => 
                           rq_vc_out_array_1_0_port, granted_vc(11) => 
                           X_Logic0_port, granted_vc(10) => 
                           granted_vc_sort_6_0_0_port, granted_vc(9) => 
                           X_Logic0_port, granted_vc(8) => X_Logic0_port, 
                           granted_vc(7) => granted_vc_sort_6_5_1_port, 
                           granted_vc(6) => granted_vc_sort_6_5_0_port, 
                           granted_vc(5) => granted_vc_sort_5_5_1_port, 
                           granted_vc(4) => granted_vc_sort_5_5_0_port, 
                           granted_vc(3) => granted_vc_sort_5_4_1_port, 
                           granted_vc(2) => granted_vc_sort_5_4_0_port, 
                           granted_vc(1) => granted_vc_sort_5_3_1_port, 
                           granted_vc(0) => granted_vc_sort_5_3_0_port, 
                           packet_end(11) => X_Logic0_port, packet_end(10) => 
                           packet_end_sort_6_0_0_port, packet_end(9) => 
                           X_Logic0_port, packet_end(8) => X_Logic0_port, 
                           packet_end(7) => packet_end_sort_6_5_1_port, 
                           packet_end(6) => packet_end_sort_6_5_0_port, 
                           packet_end(5) => packet_end_sort_5_5_1_port, 
                           packet_end(4) => packet_end_sort_5_5_0_port, 
                           packet_end(3) => packet_end_sort_5_4_1_port, 
                           packet_end(2) => packet_end_sort_5_4_0_port, 
                           packet_end(1) => packet_end_sort_5_3_1_port, 
                           packet_end(0) => packet_end_sort_5_3_0_port, 
                           crossbar_ctrl_vec(5) => crossbar_ctrl_vec(8), 
                           crossbar_ctrl_vec(4) => crossbar_ctrl_vec(7), 
                           crossbar_ctrl_vec(3) => crossbar_ctrl_vec(6), 
                           crossbar_ctrl_vec(2) => crossbar_ctrl_vec(5), 
                           crossbar_ctrl_vec(1) => crossbar_ctrl_vec(4), 
                           crossbar_ctrl_vec(0) => crossbar_ctrl_vec(3), 
                           vc_sel_enc(1) => vc_sel_enc_vec(2), vc_sel_enc(0) =>
                           vc_sel_enc_vec(1), output_vc_in_use(1) => 
                           output_vc_in_use(2), output_vc_in_use(0) => 
                           output_vc_in_use(1), ack_rq_vc_out(5) => 
                           ack_rq_vc_out_1_5_port, ack_rq_vc_out(4) => n_1763, 
                           ack_rq_vc_out(3) => ack_rq_vc_out_1_3_port, 
                           ack_rq_vc_out(2) => ack_rq_vc_out_1_2_port, 
                           ack_rq_vc_out(1) => ack_rq_vc_out_1_1_port, 
                           ack_rq_vc_out(0) => ack_rq_vc_out_1_0_port);
   input_first_arbiter_i_2 : header_arbiter_and_decoder_1_1_1_7_2_2_1_DXYU port
                           map( clk => clk, rst => n3, header(19) => header(49)
                           , header(18) => header(48), header(17) => header(47)
                           , header(16) => header(46), header(15) => header(45)
                           , header(14) => header(44), header(13) => header(43)
                           , header(12) => header(42), header(11) => header(41)
                           , header(10) => header(40), header(9) => header(39),
                           header(8) => header(38), header(7) => header(37), 
                           header(6) => header(36), header(5) => header(35), 
                           header(4) => header(34), header(3) => header(33), 
                           header(2) => header(32), header(1) => header(31), 
                           header(0) => header(30), valid_data_vc(1) => 
                           valid_data_vc_vec(4), valid_data_vc(0) => 
                           valid_data_vc_vec(3), enr_vc(1) => enr_vc(4), 
                           enr_vc(0) => enr_vc(3), ack_vc => 
                           ack_rq_vc_out_var_2_port, granted_rq(6) => n_1764, 
                           granted_rq(5) => rq_vc_out_array_5_3_port, 
                           granted_rq(4) => rq_vc_out_array_4_4_port, 
                           granted_rq(3) => rq_vc_out_array_3_5_port, 
                           granted_rq(2) => n_1765, granted_rq(1) => 
                           rq_vc_out_array_1_0_port, granted_rq(0) => 
                           rq_vc_out_array_0_1_port, input_vc_in_use(1) => 
                           input_vc_in_use(4), input_vc_in_use(0) => 
                           input_vc_in_use(3), packet_end(1) => 
                           packet_end_sort_5_3_1_port, packet_end(0) => 
                           packet_end_sort_5_3_0_port, granted_vc(1) => 
                           granted_vc_sort_5_3_1_port, granted_vc(0) => 
                           granted_vc_sort_5_3_0_port);
   output_last_arbiter_i_2 : vc_output_allocator_port_num7_vc_num_out2_5 port 
                           map( clk => clk, rst => n3, rq_vc_out(5) => 
                           X_Logic0_port, rq_vc_out(4) => 
                           rq_vc_out_array_2_4_port, rq_vc_out(3) => 
                           X_Logic0_port, rq_vc_out(2) => 
                           rq_vc_out_array_2_2_port, rq_vc_out(1) => 
                           rq_vc_out_array_2_1_port, rq_vc_out(0) => 
                           X_Logic0_port, granted_vc(11) => X_Logic0_port, 
                           granted_vc(10) => X_Logic0_port, granted_vc(9) => 
                           X_Logic0_port, granted_vc(8) => 
                           granted_vc_sort_6_0_0_port, granted_vc(7) => 
                           X_Logic0_port, granted_vc(6) => X_Logic0_port, 
                           granted_vc(5) => granted_vc_sort_6_5_1_port, 
                           granted_vc(4) => granted_vc_sort_6_5_0_port, 
                           granted_vc(3) => granted_vc_sort_5_5_1_port, 
                           granted_vc(2) => granted_vc_sort_5_5_0_port, 
                           granted_vc(1) => X_Logic0_port, granted_vc(0) => 
                           X_Logic0_port, packet_end(11) => X_Logic0_port, 
                           packet_end(10) => X_Logic0_port, packet_end(9) => 
                           X_Logic0_port, packet_end(8) => 
                           packet_end_sort_6_0_0_port, packet_end(7) => 
                           X_Logic0_port, packet_end(6) => X_Logic0_port, 
                           packet_end(5) => packet_end_sort_6_5_1_port, 
                           packet_end(4) => packet_end_sort_6_5_0_port, 
                           packet_end(3) => packet_end_sort_5_5_1_port, 
                           packet_end(2) => packet_end_sort_5_5_0_port, 
                           packet_end(1) => X_Logic0_port, packet_end(0) => 
                           X_Logic0_port, crossbar_ctrl_vec(5) => 
                           crossbar_ctrl_vec(14), crossbar_ctrl_vec(4) => 
                           crossbar_ctrl_vec(13), crossbar_ctrl_vec(3) => 
                           crossbar_ctrl_vec(12), crossbar_ctrl_vec(2) => 
                           crossbar_ctrl_vec(11), crossbar_ctrl_vec(1) => 
                           crossbar_ctrl_vec(10), crossbar_ctrl_vec(0) => 
                           crossbar_ctrl_vec(9), vc_sel_enc(1) => 
                           vc_sel_enc_vec(4), vc_sel_enc(0) => 
                           vc_sel_enc_vec(3), output_vc_in_use(1) => 
                           output_vc_in_use(4), output_vc_in_use(0) => 
                           output_vc_in_use(3), ack_rq_vc_out(5) => n_1766, 
                           ack_rq_vc_out(4) => ack_rq_vc_out_2_4_port, 
                           ack_rq_vc_out(3) => n_1767, ack_rq_vc_out(2) => 
                           ack_rq_vc_out_2_2_port, ack_rq_vc_out(1) => 
                           ack_rq_vc_out_2_1_port, ack_rq_vc_out(0) => n_1768);
   input_first_arbiter_i_3 : header_arbiter_and_decoder_1_1_1_7_3_2_1_DXYU port
                           map( clk => clk, rst => n3, header(19) => header(69)
                           , header(18) => header(68), header(17) => header(67)
                           , header(16) => header(66), header(15) => header(65)
                           , header(14) => header(64), header(13) => header(63)
                           , header(12) => header(62), header(11) => header(61)
                           , header(10) => header(60), header(9) => header(59),
                           header(8) => header(58), header(7) => header(57), 
                           header(6) => header(56), header(5) => header(55), 
                           header(4) => header(54), header(3) => header(53), 
                           header(2) => header(52), header(1) => header(51), 
                           header(0) => header(50), valid_data_vc(1) => 
                           valid_data_vc_vec(6), valid_data_vc(0) => 
                           valid_data_vc_vec(5), enr_vc(1) => enr_vc(6), 
                           enr_vc(0) => enr_vc(5), ack_vc => 
                           ack_rq_vc_out_var_3_port, granted_rq(6) => n_1769, 
                           granted_rq(5) => rq_vc_out_array_5_4_port, 
                           granted_rq(4) => n_1770, granted_rq(3) => n_1771, 
                           granted_rq(2) => n_1772, granted_rq(1) => 
                           rq_vc_out_array_1_1_port, granted_rq(0) => 
                           rq_vc_out_array_0_2_port, input_vc_in_use(1) => 
                           input_vc_in_use(6), input_vc_in_use(0) => 
                           input_vc_in_use(5), packet_end(1) => 
                           packet_end_sort_5_4_1_port, packet_end(0) => 
                           packet_end_sort_5_4_0_port, granted_vc(1) => 
                           granted_vc_sort_5_4_1_port, granted_vc(0) => 
                           granted_vc_sort_5_4_0_port);
   output_last_arbiter_i_3 : vc_output_allocator_port_num7_vc_num_out2_4 port 
                           map( clk => clk, rst => n3, rq_vc_out(5) => 
                           rq_vc_out_array_3_5_port, rq_vc_out(4) => 
                           rq_vc_out_array_3_4_port, rq_vc_out(3) => 
                           rq_vc_out_array_3_3_port, rq_vc_out(2) => 
                           X_Logic0_port, rq_vc_out(1) => 
                           rq_vc_out_array_3_1_port, rq_vc_out(0) => 
                           rq_vc_out_array_3_0_port, granted_vc(11) => 
                           granted_vc_sort_5_3_1_port, granted_vc(10) => 
                           granted_vc_sort_5_3_0_port, granted_vc(9) => 
                           granted_vc_sort_5_2_1_port, granted_vc(8) => 
                           granted_vc_sort_5_2_0_port, granted_vc(7) => 
                           X_Logic0_port, granted_vc(6) => 
                           granted_vc_sort_6_0_0_port, granted_vc(5) => 
                           X_Logic0_port, granted_vc(4) => X_Logic0_port, 
                           granted_vc(3) => granted_vc_sort_6_5_1_port, 
                           granted_vc(2) => granted_vc_sort_6_5_0_port, 
                           granted_vc(1) => granted_vc_sort_5_5_1_port, 
                           granted_vc(0) => granted_vc_sort_5_5_0_port, 
                           packet_end(11) => packet_end_sort_5_3_1_port, 
                           packet_end(10) => packet_end_sort_5_3_0_port, 
                           packet_end(9) => packet_end_sort_5_2_1_port, 
                           packet_end(8) => packet_end_sort_5_2_0_port, 
                           packet_end(7) => X_Logic0_port, packet_end(6) => 
                           packet_end_sort_6_0_0_port, packet_end(5) => 
                           X_Logic0_port, packet_end(4) => X_Logic0_port, 
                           packet_end(3) => packet_end_sort_6_5_1_port, 
                           packet_end(2) => packet_end_sort_6_5_0_port, 
                           packet_end(1) => packet_end_sort_5_5_1_port, 
                           packet_end(0) => packet_end_sort_5_5_0_port, 
                           crossbar_ctrl_vec(5) => crossbar_ctrl_vec(20), 
                           crossbar_ctrl_vec(4) => crossbar_ctrl_vec(19), 
                           crossbar_ctrl_vec(3) => crossbar_ctrl_vec(18), 
                           crossbar_ctrl_vec(2) => crossbar_ctrl_vec(17), 
                           crossbar_ctrl_vec(1) => crossbar_ctrl_vec(16), 
                           crossbar_ctrl_vec(0) => crossbar_ctrl_vec(15), 
                           vc_sel_enc(1) => vc_sel_enc_vec(6), vc_sel_enc(0) =>
                           vc_sel_enc_vec(5), output_vc_in_use(1) => 
                           output_vc_in_use(6), output_vc_in_use(0) => 
                           output_vc_in_use(5), ack_rq_vc_out(5) => 
                           ack_rq_vc_out_3_5_port, ack_rq_vc_out(4) => 
                           ack_rq_vc_out_3_4_port, ack_rq_vc_out(3) => 
                           ack_rq_vc_out_3_3_port, ack_rq_vc_out(2) => n_1773, 
                           ack_rq_vc_out(1) => ack_rq_vc_out_3_1_port, 
                           ack_rq_vc_out(0) => ack_rq_vc_out_3_0_port);
   input_first_arbiter_i_4 : header_arbiter_and_decoder_1_1_1_7_4_2_1_DXYU port
                           map( clk => clk, rst => n3, header(19) => header(89)
                           , header(18) => header(88), header(17) => header(87)
                           , header(16) => header(86), header(15) => header(85)
                           , header(14) => header(84), header(13) => header(83)
                           , header(12) => header(82), header(11) => header(81)
                           , header(10) => header(80), header(9) => header(79),
                           header(8) => header(78), header(7) => header(77), 
                           header(6) => header(76), header(5) => header(75), 
                           header(4) => header(74), header(3) => header(73), 
                           header(2) => header(72), header(1) => header(71), 
                           header(0) => header(70), valid_data_vc(1) => 
                           valid_data_vc_vec(8), valid_data_vc(0) => 
                           valid_data_vc_vec(7), enr_vc(1) => enr_vc(8), 
                           enr_vc(0) => enr_vc(7), ack_vc => 
                           ack_rq_vc_out_var_4_port, granted_rq(6) => n_1774, 
                           granted_rq(5) => rq_vc_out_array_5_5_port, 
                           granted_rq(4) => n_1775, granted_rq(3) => 
                           rq_vc_out_array_3_0_port, granted_rq(2) => 
                           rq_vc_out_array_2_1_port, granted_rq(1) => 
                           rq_vc_out_array_1_2_port, granted_rq(0) => 
                           rq_vc_out_array_0_3_port, input_vc_in_use(1) => 
                           input_vc_in_use(8), input_vc_in_use(0) => 
                           input_vc_in_use(7), packet_end(1) => 
                           packet_end_sort_5_5_1_port, packet_end(0) => 
                           packet_end_sort_5_5_0_port, granted_vc(1) => 
                           granted_vc_sort_5_5_1_port, granted_vc(0) => 
                           granted_vc_sort_5_5_0_port);
   output_last_arbiter_i_4 : vc_output_allocator_port_num7_vc_num_out2_3 port 
                           map( clk => clk, rst => n3, rq_vc_out(5) => 
                           X_Logic0_port, rq_vc_out(4) => 
                           rq_vc_out_array_4_4_port, rq_vc_out(3) => 
                           X_Logic0_port, rq_vc_out(2) => 
                           rq_vc_out_array_4_2_port, rq_vc_out(1) => 
                           X_Logic0_port, rq_vc_out(0) => 
                           rq_vc_out_array_4_0_port, granted_vc(11) => 
                           X_Logic0_port, granted_vc(10) => X_Logic0_port, 
                           granted_vc(9) => granted_vc_sort_5_3_1_port, 
                           granted_vc(8) => granted_vc_sort_5_3_0_port, 
                           granted_vc(7) => X_Logic0_port, granted_vc(6) => 
                           X_Logic0_port, granted_vc(5) => X_Logic0_port, 
                           granted_vc(4) => granted_vc_sort_6_0_0_port, 
                           granted_vc(3) => X_Logic0_port, granted_vc(2) => 
                           X_Logic0_port, granted_vc(1) => 
                           granted_vc_sort_6_5_1_port, granted_vc(0) => 
                           granted_vc_sort_6_5_0_port, packet_end(11) => 
                           X_Logic0_port, packet_end(10) => X_Logic0_port, 
                           packet_end(9) => packet_end_sort_5_3_1_port, 
                           packet_end(8) => packet_end_sort_5_3_0_port, 
                           packet_end(7) => X_Logic0_port, packet_end(6) => 
                           X_Logic0_port, packet_end(5) => X_Logic0_port, 
                           packet_end(4) => packet_end_sort_6_0_0_port, 
                           packet_end(3) => X_Logic0_port, packet_end(2) => 
                           X_Logic0_port, packet_end(1) => 
                           packet_end_sort_6_5_1_port, packet_end(0) => 
                           packet_end_sort_6_5_0_port, crossbar_ctrl_vec(5) => 
                           crossbar_ctrl_vec(26), crossbar_ctrl_vec(4) => 
                           crossbar_ctrl_vec(25), crossbar_ctrl_vec(3) => 
                           crossbar_ctrl_vec(24), crossbar_ctrl_vec(2) => 
                           crossbar_ctrl_vec(23), crossbar_ctrl_vec(1) => 
                           crossbar_ctrl_vec(22), crossbar_ctrl_vec(0) => 
                           crossbar_ctrl_vec(21), vc_sel_enc(1) => 
                           vc_sel_enc_vec(8), vc_sel_enc(0) => 
                           vc_sel_enc_vec(7), output_vc_in_use(1) => 
                           output_vc_in_use(8), output_vc_in_use(0) => 
                           output_vc_in_use(7), ack_rq_vc_out(5) => n_1776, 
                           ack_rq_vc_out(4) => ack_rq_vc_out_4_4_port, 
                           ack_rq_vc_out(3) => n_1777, ack_rq_vc_out(2) => 
                           ack_rq_vc_out_4_2_port, ack_rq_vc_out(1) => n_1778, 
                           ack_rq_vc_out(0) => ack_rq_vc_out_4_0_port);
   input_first_arbiter_i_5 : header_arbiter_and_decoder_1_1_1_7_5_2_1_DXYU port
                           map( clk => clk, rst => n3, header(19) => 
                           header(109), header(18) => header(108), header(17) 
                           => header(107), header(16) => header(106), 
                           header(15) => header(105), header(14) => header(104)
                           , header(13) => header(103), header(12) => 
                           header(102), header(11) => header(101), header(10) 
                           => header(100), header(9) => header(99), header(8) 
                           => header(98), header(7) => header(97), header(6) =>
                           header(96), header(5) => header(95), header(4) => 
                           header(94), header(3) => header(93), header(2) => 
                           header(92), header(1) => header(91), header(0) => 
                           header(90), valid_data_vc(1) => 
                           valid_data_vc_vec(10), valid_data_vc(0) => 
                           valid_data_vc_vec(9), enr_vc(1) => enr_vc(10), 
                           enr_vc(0) => enr_vc(9), ack_vc => 
                           ack_rq_vc_out_var_5_port, granted_rq(6) => 
                           rq_vc_out_array_6_5_port, granted_rq(5) => n_1779, 
                           granted_rq(4) => rq_vc_out_array_4_0_port, 
                           granted_rq(3) => rq_vc_out_array_3_1_port, 
                           granted_rq(2) => rq_vc_out_array_2_2_port, 
                           granted_rq(1) => rq_vc_out_array_1_3_port, 
                           granted_rq(0) => rq_vc_out_array_0_4_port, 
                           input_vc_in_use(1) => input_vc_in_use(10), 
                           input_vc_in_use(0) => input_vc_in_use(9), 
                           packet_end(1) => packet_end_sort_6_5_1_port, 
                           packet_end(0) => packet_end_sort_6_5_0_port, 
                           granted_vc(1) => granted_vc_sort_6_5_1_port, 
                           granted_vc(0) => granted_vc_sort_6_5_0_port);
   output_last_arbiter_i_5 : vc_output_allocator_port_num7_vc_num_out2_2 port 
                           map( clk => clk, rst => n3, rq_vc_out(5) => 
                           rq_vc_out_array_5_5_port, rq_vc_out(4) => 
                           rq_vc_out_array_5_4_port, rq_vc_out(3) => 
                           rq_vc_out_array_5_3_port, rq_vc_out(2) => 
                           rq_vc_out_array_5_2_port, rq_vc_out(1) => 
                           rq_vc_out_array_5_1_port, rq_vc_out(0) => 
                           rq_vc_out_array_5_0_port, granted_vc(11) => 
                           granted_vc_sort_5_5_1_port, granted_vc(10) => 
                           granted_vc_sort_5_5_0_port, granted_vc(9) => 
                           granted_vc_sort_5_4_1_port, granted_vc(8) => 
                           granted_vc_sort_5_4_0_port, granted_vc(7) => 
                           granted_vc_sort_5_3_1_port, granted_vc(6) => 
                           granted_vc_sort_5_3_0_port, granted_vc(5) => 
                           granted_vc_sort_5_2_1_port, granted_vc(4) => 
                           granted_vc_sort_5_2_0_port, granted_vc(3) => 
                           X_Logic0_port, granted_vc(2) => 
                           granted_vc_sort_6_0_0_port, granted_vc(1) => 
                           granted_vc_sort_5_0_1_port, granted_vc(0) => 
                           granted_vc_sort_5_0_0_port, packet_end(11) => 
                           packet_end_sort_5_5_1_port, packet_end(10) => 
                           packet_end_sort_5_5_0_port, packet_end(9) => 
                           packet_end_sort_5_4_1_port, packet_end(8) => 
                           packet_end_sort_5_4_0_port, packet_end(7) => 
                           packet_end_sort_5_3_1_port, packet_end(6) => 
                           packet_end_sort_5_3_0_port, packet_end(5) => 
                           packet_end_sort_5_2_1_port, packet_end(4) => 
                           packet_end_sort_5_2_0_port, packet_end(3) => 
                           X_Logic0_port, packet_end(2) => 
                           packet_end_sort_6_0_0_port, packet_end(1) => 
                           packet_end_sort_5_0_1_port, packet_end(0) => 
                           packet_end_sort_5_0_0_port, crossbar_ctrl_vec(5) => 
                           crossbar_ctrl_vec(32), crossbar_ctrl_vec(4) => 
                           crossbar_ctrl_vec(31), crossbar_ctrl_vec(3) => 
                           crossbar_ctrl_vec(30), crossbar_ctrl_vec(2) => 
                           crossbar_ctrl_vec(29), crossbar_ctrl_vec(1) => 
                           crossbar_ctrl_vec(28), crossbar_ctrl_vec(0) => 
                           crossbar_ctrl_vec(27), vc_sel_enc(1) => 
                           vc_sel_enc_vec(10), vc_sel_enc(0) => 
                           vc_sel_enc_vec(9), output_vc_in_use(1) => 
                           output_vc_in_use(10), output_vc_in_use(0) => 
                           output_vc_in_use(9), ack_rq_vc_out(5) => 
                           ack_rq_vc_out_5_5_port, ack_rq_vc_out(4) => 
                           ack_rq_vc_out_5_4_port, ack_rq_vc_out(3) => 
                           ack_rq_vc_out_5_3_port, ack_rq_vc_out(2) => 
                           ack_rq_vc_out_5_2_port, ack_rq_vc_out(1) => 
                           ack_rq_vc_out_5_1_port, ack_rq_vc_out(0) => 
                           ack_rq_vc_out_5_0_port);
   input_first_arbiter_i_6 : header_arbiter_and_decoder_1_1_1_7_6_2_1_DXYU port
                           map( clk => clk, rst => n3, header(19) => 
                           header(129), header(18) => header(128), header(17) 
                           => header(127), header(16) => header(126), 
                           header(15) => header(125), header(14) => header(124)
                           , header(13) => header(123), header(12) => 
                           header(122), header(11) => header(121), header(10) 
                           => header(120), header(9) => header(119), header(8) 
                           => header(118), header(7) => header(117), header(6) 
                           => header(116), header(5) => header(115), header(4) 
                           => header(114), header(3) => header(113), header(2) 
                           => header(112), header(1) => header(111), header(0) 
                           => header(110), valid_data_vc(1) => 
                           valid_data_vc_vec(12), valid_data_vc(0) => 
                           valid_data_vc_vec(11), enr_vc(1) => enr_vc(12), 
                           enr_vc(0) => enr_vc(11), ack_vc => 
                           ack_rq_vc_out_var_6_port, granted_rq(6) => n_1780, 
                           granted_rq(5) => rq_vc_out_array_5_0_port, 
                           granted_rq(4) => n_1781, granted_rq(3) => n_1782, 
                           granted_rq(2) => n_1783, granted_rq(1) => n_1784, 
                           granted_rq(0) => rq_vc_out_array_0_5_port, 
                           input_vc_in_use(1) => input_vc_in_use(12), 
                           input_vc_in_use(0) => input_vc_in_use(11), 
                           packet_end(1) => packet_end_sort_5_0_1_port, 
                           packet_end(0) => packet_end_sort_5_0_0_port, 
                           granted_vc(1) => granted_vc_sort_5_0_1_port, 
                           granted_vc(0) => granted_vc_sort_5_0_0_port);
   output_last_arbiter_i_6 : vc_output_allocator_port_num7_vc_num_out2_1 port 
                           map( clk => clk, rst => n3, rq_vc_out(5) => 
                           rq_vc_out_array_6_5_port, rq_vc_out(4) => 
                           X_Logic0_port, rq_vc_out(3) => X_Logic0_port, 
                           rq_vc_out(2) => X_Logic0_port, rq_vc_out(1) => 
                           X_Logic0_port, rq_vc_out(0) => 
                           rq_vc_out_array_6_0_port, granted_vc(11) => 
                           granted_vc_sort_6_5_1_port, granted_vc(10) => 
                           granted_vc_sort_6_5_0_port, granted_vc(9) => 
                           X_Logic0_port, granted_vc(8) => X_Logic0_port, 
                           granted_vc(7) => X_Logic0_port, granted_vc(6) => 
                           X_Logic0_port, granted_vc(5) => X_Logic0_port, 
                           granted_vc(4) => X_Logic0_port, granted_vc(3) => 
                           X_Logic0_port, granted_vc(2) => X_Logic0_port, 
                           granted_vc(1) => X_Logic0_port, granted_vc(0) => 
                           granted_vc_sort_6_0_0_port, packet_end(11) => 
                           packet_end_sort_6_5_1_port, packet_end(10) => 
                           packet_end_sort_6_5_0_port, packet_end(9) => 
                           X_Logic0_port, packet_end(8) => X_Logic0_port, 
                           packet_end(7) => X_Logic0_port, packet_end(6) => 
                           X_Logic0_port, packet_end(5) => X_Logic0_port, 
                           packet_end(4) => X_Logic0_port, packet_end(3) => 
                           X_Logic0_port, packet_end(2) => X_Logic0_port, 
                           packet_end(1) => X_Logic0_port, packet_end(0) => 
                           packet_end_sort_6_0_0_port, crossbar_ctrl_vec(5) => 
                           crossbar_ctrl_vec(38), crossbar_ctrl_vec(4) => 
                           crossbar_ctrl_vec(37), crossbar_ctrl_vec(3) => 
                           crossbar_ctrl_vec(36), crossbar_ctrl_vec(2) => 
                           crossbar_ctrl_vec(35), crossbar_ctrl_vec(1) => 
                           crossbar_ctrl_vec(34), crossbar_ctrl_vec(0) => 
                           crossbar_ctrl_vec(33), vc_sel_enc(1) => 
                           vc_sel_enc_vec(12), vc_sel_enc(0) => 
                           vc_sel_enc_vec(11), output_vc_in_use(1) => 
                           output_vc_in_use(12), output_vc_in_use(0) => 
                           output_vc_in_use(11), ack_rq_vc_out(5) => 
                           ack_rq_vc_out_6_5_port, ack_rq_vc_out(4) => n_1785, 
                           ack_rq_vc_out(3) => n_1786, ack_rq_vc_out(2) => 
                           n_1787, ack_rq_vc_out(1) => n_1788, ack_rq_vc_out(0)
                           => ack_rq_vc_out_6_0_port);
   U11 : HB1xp67_ASAP7_75t_R port map( A => rst, Y => n3);
   U12 : TIELOx1_ASAP7_75t_R port map( L => X_Logic0_port);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity fifo_buff_depth2_0 is

   port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, clk, 
         rst : in std_logic;  data_out : out std_logic_vector (63 downto 0);  
         valid_data : out std_logic);

end fifo_buff_depth2_0;

architecture SYN_rtl of fifo_buff_depth2_0 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx3_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component O2A1O1Ixp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal valid_data_port, read_pointer_0_port, fifo_1_63_port, fifo_1_62_port,
      fifo_1_61_port, fifo_1_60_port, fifo_1_59_port, fifo_1_58_port, 
      fifo_1_57_port, fifo_1_56_port, fifo_1_55_port, fifo_1_54_port, 
      fifo_1_53_port, fifo_1_52_port, fifo_1_51_port, fifo_1_50_port, 
      fifo_1_49_port, fifo_1_48_port, fifo_1_47_port, fifo_1_46_port, 
      fifo_1_45_port, fifo_1_44_port, fifo_1_43_port, fifo_1_42_port, 
      fifo_1_41_port, fifo_1_40_port, fifo_1_39_port, fifo_1_38_port, 
      fifo_1_37_port, fifo_1_36_port, fifo_1_35_port, fifo_1_34_port, 
      fifo_1_33_port, fifo_1_32_port, fifo_1_31_port, fifo_1_30_port, 
      fifo_1_29_port, fifo_1_28_port, fifo_1_27_port, fifo_1_26_port, 
      fifo_1_25_port, fifo_1_24_port, fifo_1_23_port, fifo_1_22_port, 
      fifo_1_21_port, fifo_1_20_port, fifo_1_19_port, fifo_1_18_port, 
      fifo_1_17_port, fifo_1_16_port, fifo_1_15_port, fifo_1_14_port, 
      fifo_1_13_port, fifo_1_12_port, fifo_1_11_port, fifo_1_10_port, 
      fifo_1_9_port, fifo_1_8_port, fifo_1_7_port, fifo_1_6_port, fifo_1_5_port
      , fifo_1_4_port, fifo_1_3_port, fifo_1_2_port, fifo_1_1_port, 
      fifo_1_0_port, fifo_0_63_port, fifo_0_62_port, fifo_0_61_port, 
      fifo_0_60_port, fifo_0_59_port, fifo_0_58_port, fifo_0_57_port, 
      fifo_0_56_port, fifo_0_55_port, fifo_0_54_port, fifo_0_53_port, 
      fifo_0_52_port, fifo_0_51_port, fifo_0_50_port, fifo_0_49_port, 
      fifo_0_48_port, fifo_0_47_port, fifo_0_46_port, fifo_0_45_port, 
      fifo_0_44_port, fifo_0_43_port, fifo_0_42_port, fifo_0_41_port, 
      fifo_0_40_port, fifo_0_39_port, fifo_0_38_port, fifo_0_37_port, 
      fifo_0_36_port, fifo_0_35_port, fifo_0_34_port, fifo_0_33_port, 
      fifo_0_32_port, fifo_0_31_port, fifo_0_30_port, fifo_0_29_port, 
      fifo_0_28_port, fifo_0_27_port, fifo_0_26_port, fifo_0_25_port, 
      fifo_0_24_port, fifo_0_23_port, fifo_0_22_port, fifo_0_21_port, 
      fifo_0_20_port, fifo_0_19_port, fifo_0_18_port, fifo_0_17_port, 
      fifo_0_16_port, fifo_0_15_port, fifo_0_14_port, fifo_0_13_port, 
      fifo_0_12_port, fifo_0_11_port, fifo_0_10_port, fifo_0_9_port, 
      fifo_0_8_port, fifo_0_7_port, fifo_0_6_port, fifo_0_5_port, fifo_0_4_port
      , fifo_0_3_port, fifo_0_2_port, fifo_0_1_port, fifo_0_0_port, N7, N9, n2,
      n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30, n32, 
      n34, n36, n38, n40, n42, n44, n46, n48, n50, n52, n54, n56, n58, n60, n62
      , n64, n66, n68, n70, n72, n74, n76, n78, n80, n82, n84, n86, n88, n90, 
      n92, n94, n96, n98, n100, n102, n104, n106, n108, n110, n112, n114, n116,
      n118, n120, n122, n124, n126, n128, n130, n132, n134, n136, n138, n140, 
      n142, n144, n146, n148, n150, n152, n154, n156, n158, n160, n162, n164, 
      n166, n168, n170, n172, n174, n176, n178, n180, n182, n184, n186, n188, 
      n190, n192, n194, n196, n198, n200, n202, n204, n206, n208, n210, n212, 
      n214, n216, n218, n220, n222, n224, n226, n228, n230, n232, n234, n236, 
      n238, n240, n242, n244, n246, n248, n250, n252, n254, n256, n258, n260, 
      n262, n264, n266, n268, n1, n3, n5, n7_port, n9_port, n11, n13, n15, n17,
      n19, n21, n23, n25, n27, n29, n31, n33, n35, n37, n39, n41, n43, n45, n47
      , n49 : std_logic;

begin
   valid_data <= valid_data_port;
   
   U4 : XOR2xp5_ASAP7_75t_R port map( A => N7, B => n43, Y => n2);
   U143 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_9_port, B1 => 
                           n43, B2 => fifo_0_9_port, Y => data_out(9));
   U144 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_8_port, B1 => 
                           n43, B2 => fifo_0_8_port, Y => data_out(8));
   U145 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_7_port, B1 => 
                           n43, B2 => fifo_0_7_port, Y => data_out(7));
   U146 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_6_port, B1 => 
                           n43, B2 => fifo_0_6_port, Y => data_out(6));
   U147 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_63_port, B1 => 
                           n43, B2 => fifo_0_63_port, Y => data_out(63));
   U148 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_62_port, B1 => 
                           n43, B2 => fifo_0_62_port, Y => data_out(62));
   U149 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_61_port, B1 => 
                           n43, B2 => fifo_0_61_port, Y => data_out(61));
   U150 : AO22x1_ASAP7_75t_R port map( A1 => n31, A2 => fifo_1_60_port, B1 => 
                           n43, B2 => fifo_0_60_port, Y => data_out(60));
   U151 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_5_port, B1 => 
                           n43, B2 => fifo_0_5_port, Y => data_out(5));
   U152 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_59_port, B1 => 
                           n43, B2 => fifo_0_59_port, Y => data_out(59));
   U153 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_58_port, B1 => 
                           n43, B2 => fifo_0_58_port, Y => data_out(58));
   U154 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_57_port, B1 => 
                           n43, B2 => fifo_0_57_port, Y => data_out(57));
   U155 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_56_port, B1 => 
                           n43, B2 => fifo_0_56_port, Y => data_out(56));
   U156 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_55_port, B1 => 
                           n43, B2 => fifo_0_55_port, Y => data_out(55));
   U157 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_54_port, B1 => 
                           n43, B2 => fifo_0_54_port, Y => data_out(54));
   U158 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_53_port, B1 => 
                           n43, B2 => fifo_0_53_port, Y => data_out(53));
   U159 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_52_port, B1 => 
                           n43, B2 => fifo_0_52_port, Y => data_out(52));
   U160 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_51_port, B1 => 
                           n43, B2 => fifo_0_51_port, Y => data_out(51));
   U161 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_50_port, B1 => 
                           n43, B2 => fifo_0_50_port, Y => data_out(50));
   U162 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_4_port, B1 => 
                           n43, B2 => fifo_0_4_port, Y => data_out(4));
   U163 : AO22x1_ASAP7_75t_R port map( A1 => n33, A2 => fifo_1_49_port, B1 => 
                           n43, B2 => fifo_0_49_port, Y => data_out(49));
   U164 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_48_port, B1 => 
                           n43, B2 => fifo_0_48_port, Y => data_out(48));
   U165 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_47_port, B1 => 
                           n43, B2 => fifo_0_47_port, Y => data_out(47));
   U166 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_46_port, B1 => 
                           n43, B2 => fifo_0_46_port, Y => data_out(46));
   U167 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_45_port, B1 => 
                           n43, B2 => fifo_0_45_port, Y => data_out(45));
   U168 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_44_port, B1 => 
                           n43, B2 => fifo_0_44_port, Y => data_out(44));
   U169 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_43_port, B1 => 
                           n43, B2 => fifo_0_43_port, Y => data_out(43));
   U170 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_42_port, B1 => 
                           n43, B2 => fifo_0_42_port, Y => data_out(42));
   U171 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_41_port, B1 => 
                           n43, B2 => fifo_0_41_port, Y => data_out(41));
   U172 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_40_port, B1 => 
                           n43, B2 => fifo_0_40_port, Y => data_out(40));
   U173 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_3_port, B1 => 
                           n43, B2 => fifo_0_3_port, Y => data_out(3));
   U174 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_39_port, B1 => 
                           n43, B2 => fifo_0_39_port, Y => data_out(39));
   U175 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_38_port, B1 => 
                           n43, B2 => fifo_0_38_port, Y => data_out(38));
   U176 : AO22x1_ASAP7_75t_R port map( A1 => n35, A2 => fifo_1_37_port, B1 => 
                           n43, B2 => fifo_0_37_port, Y => data_out(37));
   U177 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_36_port, B1 => 
                           n43, B2 => fifo_0_36_port, Y => data_out(36));
   U178 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_35_port, B1 => 
                           n43, B2 => fifo_0_35_port, Y => data_out(35));
   U179 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_34_port, B1 => 
                           n43, B2 => fifo_0_34_port, Y => data_out(34));
   U180 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_33_port, B1 => 
                           n43, B2 => fifo_0_33_port, Y => data_out(33));
   U181 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_32_port, B1 => 
                           n43, B2 => fifo_0_32_port, Y => data_out(32));
   U182 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_31_port, B1 => 
                           n43, B2 => fifo_0_31_port, Y => data_out(31));
   U183 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_30_port, B1 => 
                           n43, B2 => fifo_0_30_port, Y => data_out(30));
   U184 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_2_port, B1 => 
                           n43, B2 => fifo_0_2_port, Y => data_out(2));
   U185 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_29_port, B1 => 
                           n43, B2 => fifo_0_29_port, Y => data_out(29));
   U186 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_28_port, B1 => 
                           n43, B2 => fifo_0_28_port, Y => data_out(28));
   U187 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_27_port, B1 => 
                           n43, B2 => fifo_0_27_port, Y => data_out(27));
   U188 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_26_port, B1 => 
                           n43, B2 => fifo_0_26_port, Y => data_out(26));
   U189 : AO22x1_ASAP7_75t_R port map( A1 => n37, A2 => fifo_1_25_port, B1 => 
                           n43, B2 => fifo_0_25_port, Y => data_out(25));
   U190 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_24_port, B1 => 
                           n43, B2 => fifo_0_24_port, Y => data_out(24));
   U191 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_23_port, B1 => 
                           n43, B2 => fifo_0_23_port, Y => data_out(23));
   U192 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_22_port, B1 => 
                           n43, B2 => fifo_0_22_port, Y => data_out(22));
   U193 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_21_port, B1 => 
                           n43, B2 => fifo_0_21_port, Y => data_out(21));
   U194 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_20_port, B1 => 
                           n43, B2 => fifo_0_20_port, Y => data_out(20));
   U195 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_1_port, B1 => 
                           n43, B2 => fifo_0_1_port, Y => data_out(1));
   U196 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_19_port, B1 => 
                           n43, B2 => fifo_0_19_port, Y => data_out(19));
   U197 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_18_port, B1 => 
                           n43, B2 => fifo_0_18_port, Y => data_out(18));
   U198 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_17_port, B1 => 
                           n43, B2 => fifo_0_17_port, Y => data_out(17));
   U199 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_16_port, B1 => 
                           n43, B2 => fifo_0_16_port, Y => data_out(16));
   U200 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_15_port, B1 => 
                           n43, B2 => fifo_0_15_port, Y => data_out(15));
   U201 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_14_port, B1 => 
                           n43, B2 => fifo_0_14_port, Y => data_out(14));
   U202 : AO22x1_ASAP7_75t_R port map( A1 => n39, A2 => fifo_1_13_port, B1 => 
                           n43, B2 => fifo_0_13_port, Y => data_out(13));
   U203 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_12_port, B1 => 
                           n43, B2 => fifo_0_12_port, Y => data_out(12));
   U204 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_11_port, B1 => 
                           n43, B2 => fifo_0_11_port, Y => data_out(11));
   U205 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_10_port, B1 => 
                           n43, B2 => fifo_0_10_port, Y => data_out(10));
   U206 : AO22x1_ASAP7_75t_R port map( A1 => n41, A2 => fifo_1_0_port, B1 => 
                           n43, B2 => fifo_0_0_port, Y => data_out(0));
   U3 : O2A1O1Ixp5_ASAP7_75t_R port map( A1 => n47, A2 => n2, B => 
                           valid_data_port, C => write_en, Y => n8);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_0_port, A2 => n17, B1 => 
                           data_in(0), B2 => n29, Y => n10);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_1_port, A2 => n17, B1 => 
                           data_in(1), B2 => n29, Y => n12);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_2_port, A2 => n17, B1 => 
                           data_in(2), B2 => n29, Y => n14);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_3_port, A2 => n17, B1 => 
                           data_in(3), B2 => n29, Y => n16);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_4_port, A2 => n17, B1 => 
                           data_in(4), B2 => n27, Y => n18);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_5_port, A2 => n17, B1 => 
                           data_in(5), B2 => n27, Y => n20);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_6_port, A2 => n17, B1 => 
                           data_in(6), B2 => n27, Y => n22);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_7_port, A2 => n17, B1 => 
                           data_in(7), B2 => n27, Y => n24);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_8_port, A2 => n17, B1 => 
                           data_in(8), B2 => n27, Y => n26);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_9_port, A2 => n17, B1 => 
                           data_in(9), B2 => n27, Y => n28);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_10_port, A2 => n17, B1 => 
                           data_in(10), B2 => n27, Y => n30);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_11_port, A2 => n17, B1 => 
                           data_in(11), B2 => n27, Y => n32);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_12_port, A2 => n17, B1 => 
                           data_in(12), B2 => n27, Y => n34);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_13_port, A2 => n17, B1 => 
                           data_in(13), B2 => n27, Y => n36);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_14_port, A2 => n17, B1 => 
                           data_in(14), B2 => n27, Y => n38);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_15_port, A2 => n17, B1 => 
                           data_in(15), B2 => n27, Y => n40);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_16_port, A2 => n17, B1 => 
                           data_in(16), B2 => n25, Y => n42);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_17_port, A2 => n17, B1 => 
                           data_in(17), B2 => n25, Y => n44);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_18_port, A2 => n17, B1 => 
                           data_in(18), B2 => n25, Y => n46);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_19_port, A2 => n17, B1 => 
                           data_in(19), B2 => n25, Y => n48);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_20_port, A2 => n17, B1 => 
                           data_in(20), B2 => n25, Y => n50);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_21_port, A2 => n17, B1 => 
                           data_in(21), B2 => n25, Y => n52);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_22_port, A2 => n17, B1 => 
                           data_in(22), B2 => n25, Y => n54);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_23_port, A2 => n17, B1 => 
                           data_in(23), B2 => n25, Y => n56);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_24_port, A2 => n17, B1 => 
                           data_in(24), B2 => n25, Y => n58);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_25_port, A2 => n17, B1 => 
                           data_in(25), B2 => n25, Y => n60);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_26_port, A2 => n17, B1 => 
                           data_in(26), B2 => n25, Y => n62);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_27_port, A2 => n17, B1 => 
                           data_in(27), B2 => n25, Y => n64);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_28_port, A2 => n17, B1 => 
                           data_in(28), B2 => n23, Y => n66);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_29_port, A2 => n17, B1 => 
                           data_in(29), B2 => n23, Y => n68);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_30_port, A2 => n17, B1 => 
                           data_in(30), B2 => n23, Y => n70);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_31_port, A2 => n17, B1 => 
                           data_in(31), B2 => n23, Y => n72);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_32_port, A2 => n17, B1 => 
                           data_in(32), B2 => n23, Y => n74);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_33_port, A2 => n17, B1 => 
                           data_in(33), B2 => n23, Y => n76);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_34_port, A2 => n17, B1 => 
                           data_in(34), B2 => n23, Y => n78);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_35_port, A2 => n17, B1 => 
                           data_in(35), B2 => n23, Y => n80);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_36_port, A2 => n17, B1 => 
                           data_in(36), B2 => n23, Y => n82);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_37_port, A2 => n17, B1 => 
                           data_in(37), B2 => n23, Y => n84);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_38_port, A2 => n17, B1 => 
                           data_in(38), B2 => n23, Y => n86);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_39_port, A2 => n17, B1 => 
                           data_in(39), B2 => n23, Y => n88);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_40_port, A2 => n17, B1 => 
                           data_in(40), B2 => n21, Y => n90);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_41_port, A2 => n17, B1 => 
                           data_in(41), B2 => n21, Y => n92);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_42_port, A2 => n17, B1 => 
                           data_in(42), B2 => n21, Y => n94);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_43_port, A2 => n17, B1 => 
                           data_in(43), B2 => n21, Y => n96);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_44_port, A2 => n17, B1 => 
                           data_in(44), B2 => n21, Y => n98);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_45_port, A2 => n17, B1 => 
                           data_in(45), B2 => n21, Y => n100);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_46_port, A2 => n17, B1 => 
                           data_in(46), B2 => n21, Y => n102);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_47_port, A2 => n17, B1 => 
                           data_in(47), B2 => n21, Y => n104);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_48_port, A2 => n17, B1 => 
                           data_in(48), B2 => n21, Y => n106);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_49_port, A2 => n17, B1 => 
                           data_in(49), B2 => n21, Y => n108);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_50_port, A2 => n17, B1 => 
                           data_in(50), B2 => n21, Y => n110);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_51_port, A2 => n17, B1 => 
                           data_in(51), B2 => n21, Y => n112);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_52_port, A2 => n17, B1 => 
                           data_in(52), B2 => n19, Y => n114);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_53_port, A2 => n17, B1 => 
                           data_in(53), B2 => n19, Y => n116);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_54_port, A2 => n17, B1 => 
                           data_in(54), B2 => n19, Y => n118);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_55_port, A2 => n17, B1 => 
                           data_in(55), B2 => n19, Y => n120);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_56_port, A2 => n17, B1 => 
                           data_in(56), B2 => n19, Y => n122);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_57_port, A2 => n17, B1 => 
                           data_in(57), B2 => n19, Y => n124);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_58_port, A2 => n17, B1 => 
                           data_in(58), B2 => n19, Y => n126);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_59_port, A2 => n17, B1 => 
                           data_in(59), B2 => n19, Y => n128);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_60_port, A2 => n17, B1 => 
                           data_in(60), B2 => n19, Y => n130);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_61_port, A2 => n17, B1 => 
                           data_in(61), B2 => n19, Y => n132);
   U67 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_62_port, A2 => n17, B1 => 
                           data_in(62), B2 => n19, Y => n134);
   U68 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_0_63_port, A2 => n17, B1 => 
                           data_in(63), B2 => n19, Y => n136);
   U70 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N9, Y => n4);
   U71 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_0_port, A2 => n3, B1 => 
                           data_in(0), B2 => n15, Y => n138);
   U72 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_1_port, A2 => n3, B1 => 
                           data_in(1), B2 => n15, Y => n140);
   U73 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_2_port, A2 => n3, B1 => 
                           data_in(2), B2 => n15, Y => n142);
   U74 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_3_port, A2 => n3, B1 => 
                           data_in(3), B2 => n15, Y => n144);
   U75 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_4_port, A2 => n3, B1 => 
                           data_in(4), B2 => n13, Y => n146);
   U76 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_5_port, A2 => n3, B1 => 
                           data_in(5), B2 => n13, Y => n148);
   U77 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_6_port, A2 => n3, B1 => 
                           data_in(6), B2 => n13, Y => n150);
   U78 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_7_port, A2 => n3, B1 => 
                           data_in(7), B2 => n13, Y => n152);
   U79 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_8_port, A2 => n3, B1 => 
                           data_in(8), B2 => n13, Y => n154);
   U80 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_9_port, A2 => n3, B1 => 
                           data_in(9), B2 => n13, Y => n156);
   U81 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_10_port, A2 => n3, B1 => 
                           data_in(10), B2 => n13, Y => n158);
   U82 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_11_port, A2 => n3, B1 => 
                           data_in(11), B2 => n13, Y => n160);
   U83 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_12_port, A2 => n3, B1 => 
                           data_in(12), B2 => n13, Y => n162);
   U84 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_13_port, A2 => n3, B1 => 
                           data_in(13), B2 => n13, Y => n164);
   U85 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_14_port, A2 => n3, B1 => 
                           data_in(14), B2 => n13, Y => n166);
   U86 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_15_port, A2 => n3, B1 => 
                           data_in(15), B2 => n13, Y => n168);
   U87 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_16_port, A2 => n3, B1 => 
                           data_in(16), B2 => n11, Y => n170);
   U88 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_17_port, A2 => n3, B1 => 
                           data_in(17), B2 => n11, Y => n172);
   U89 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_18_port, A2 => n3, B1 => 
                           data_in(18), B2 => n11, Y => n174);
   U90 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_19_port, A2 => n3, B1 => 
                           data_in(19), B2 => n11, Y => n176);
   U91 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_20_port, A2 => n3, B1 => 
                           data_in(20), B2 => n11, Y => n178);
   U92 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_21_port, A2 => n3, B1 => 
                           data_in(21), B2 => n11, Y => n180);
   U93 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_22_port, A2 => n3, B1 => 
                           data_in(22), B2 => n11, Y => n182);
   U94 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_23_port, A2 => n3, B1 => 
                           data_in(23), B2 => n11, Y => n184);
   U95 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_24_port, A2 => n3, B1 => 
                           data_in(24), B2 => n11, Y => n186);
   U96 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_25_port, A2 => n3, B1 => 
                           data_in(25), B2 => n11, Y => n188);
   U97 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_26_port, A2 => n3, B1 => 
                           data_in(26), B2 => n11, Y => n190);
   U98 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_27_port, A2 => n3, B1 => 
                           data_in(27), B2 => n11, Y => n192);
   U99 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_28_port, A2 => n3, B1 => 
                           data_in(28), B2 => n9_port, Y => n194);
   U100 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_29_port, A2 => n3, B1 => 
                           data_in(29), B2 => n9_port, Y => n196);
   U101 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_30_port, A2 => n3, B1 => 
                           data_in(30), B2 => n9_port, Y => n198);
   U102 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_31_port, A2 => n3, B1 => 
                           data_in(31), B2 => n9_port, Y => n200);
   U103 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_32_port, A2 => n3, B1 => 
                           data_in(32), B2 => n9_port, Y => n202);
   U104 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_33_port, A2 => n3, B1 => 
                           data_in(33), B2 => n9_port, Y => n204);
   U105 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_34_port, A2 => n3, B1 => 
                           data_in(34), B2 => n9_port, Y => n206);
   U106 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_35_port, A2 => n3, B1 => 
                           data_in(35), B2 => n9_port, Y => n208);
   U107 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_36_port, A2 => n3, B1 => 
                           data_in(36), B2 => n9_port, Y => n210);
   U108 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_37_port, A2 => n3, B1 => 
                           data_in(37), B2 => n9_port, Y => n212);
   U109 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_38_port, A2 => n3, B1 => 
                           data_in(38), B2 => n9_port, Y => n214);
   U110 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_39_port, A2 => n3, B1 => 
                           data_in(39), B2 => n9_port, Y => n216);
   U111 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_40_port, A2 => n3, B1 => 
                           data_in(40), B2 => n7_port, Y => n218);
   U112 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_41_port, A2 => n3, B1 => 
                           data_in(41), B2 => n7_port, Y => n220);
   U113 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_42_port, A2 => n3, B1 => 
                           data_in(42), B2 => n7_port, Y => n222);
   U114 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_43_port, A2 => n3, B1 => 
                           data_in(43), B2 => n7_port, Y => n224);
   U115 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_44_port, A2 => n3, B1 => 
                           data_in(44), B2 => n7_port, Y => n226);
   U116 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_45_port, A2 => n3, B1 => 
                           data_in(45), B2 => n7_port, Y => n228);
   U117 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_46_port, A2 => n3, B1 => 
                           data_in(46), B2 => n7_port, Y => n230);
   U118 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_47_port, A2 => n3, B1 => 
                           data_in(47), B2 => n7_port, Y => n232);
   U119 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_48_port, A2 => n3, B1 => 
                           data_in(48), B2 => n7_port, Y => n234);
   U120 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_49_port, A2 => n3, B1 => 
                           data_in(49), B2 => n7_port, Y => n236);
   U121 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_50_port, A2 => n3, B1 => 
                           data_in(50), B2 => n7_port, Y => n238);
   U122 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_51_port, A2 => n3, B1 => 
                           data_in(51), B2 => n7_port, Y => n240);
   U123 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_52_port, A2 => n3, B1 => 
                           data_in(52), B2 => n5, Y => n242);
   U124 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_53_port, A2 => n3, B1 => 
                           data_in(53), B2 => n5, Y => n244);
   U125 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_54_port, A2 => n3, B1 => 
                           data_in(54), B2 => n5, Y => n246);
   U126 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_55_port, A2 => n3, B1 => 
                           data_in(55), B2 => n5, Y => n248);
   U127 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_56_port, A2 => n3, B1 => 
                           data_in(56), B2 => n5, Y => n250);
   U128 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_57_port, A2 => n3, B1 => 
                           data_in(57), B2 => n5, Y => n252);
   U129 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_58_port, A2 => n3, B1 => 
                           data_in(58), B2 => n5, Y => n254);
   U130 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_59_port, A2 => n3, B1 => 
                           data_in(59), B2 => n5, Y => n256);
   U131 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_60_port, A2 => n3, B1 => 
                           data_in(60), B2 => n5, Y => n258);
   U132 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_61_port, A2 => n3, B1 => 
                           data_in(61), B2 => n5, Y => n260);
   U133 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_62_port, A2 => n3, B1 => 
                           data_in(62), B2 => n5, Y => n262);
   U134 : OAI22xp5_ASAP7_75t_R port map( A1 => fifo_1_63_port, A2 => n3, B1 => 
                           data_in(63), B2 => n5, Y => n264);
   U136 : NAND2xp5_ASAP7_75t_R port map( A => write_en, B => N7, Y => n6);
   U137 : OAI22xp5_ASAP7_75t_R port map( A1 => n31, A2 => read_en, B1 => n43, 
                           B2 => n47, Y => n266);
   U139 : OAI22xp5_ASAP7_75t_R port map( A1 => N9, A2 => n49, B1 => write_en, 
                           B2 => N7, Y => n268);
   write_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n268, CLK
                           => clk, RESET => n45, SET => n1, QN => N7);
   fifo_reg_1_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n264, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_63_port);
   fifo_reg_1_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n262, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_62_port);
   fifo_reg_1_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n260, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_61_port);
   fifo_reg_1_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n258, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_60_port);
   fifo_reg_0_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n136, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_63_port);
   fifo_reg_0_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n134, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_62_port);
   fifo_reg_0_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n132, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_61_port);
   fifo_reg_0_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n130, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_60_port);
   fifo_reg_1_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n144, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_3_port);
   fifo_reg_1_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n142, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_2_port);
   fifo_reg_1_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n140, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_1_port);
   fifo_reg_1_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n138, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_0_port);
   fifo_reg_1_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n256, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_59_port);
   fifo_reg_1_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n254, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_58_port);
   fifo_reg_1_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n252, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_57_port);
   fifo_reg_1_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n250, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_56_port);
   fifo_reg_1_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n248, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_55_port);
   fifo_reg_1_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n246, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_54_port);
   fifo_reg_1_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n244, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_53_port);
   fifo_reg_1_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n242, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_52_port);
   fifo_reg_1_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n240, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_51_port);
   fifo_reg_1_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n238, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_50_port);
   fifo_reg_1_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n236, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_49_port);
   fifo_reg_1_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n234, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_48_port);
   fifo_reg_1_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n232, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_47_port);
   fifo_reg_1_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n230, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_46_port);
   fifo_reg_1_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n228, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_45_port);
   fifo_reg_1_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n226, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_44_port);
   fifo_reg_1_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n224, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_43_port);
   fifo_reg_1_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n222, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_42_port);
   fifo_reg_1_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n220, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_41_port);
   fifo_reg_1_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n218, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_40_port);
   fifo_reg_1_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n216, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_39_port);
   fifo_reg_1_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n214, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_38_port);
   fifo_reg_1_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n212, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_37_port);
   fifo_reg_1_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n210, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_36_port);
   fifo_reg_1_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n208, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_35_port);
   fifo_reg_1_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n206, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_34_port);
   fifo_reg_1_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n204, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_33_port);
   fifo_reg_1_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n202, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_32_port);
   fifo_reg_1_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n200, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_31_port);
   fifo_reg_1_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n198, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_30_port);
   fifo_reg_1_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n196, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_29_port);
   fifo_reg_1_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n194, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_28_port);
   fifo_reg_1_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n192, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_27_port);
   fifo_reg_1_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n190, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_26_port);
   fifo_reg_1_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n188, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_25_port);
   fifo_reg_1_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n186, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_24_port);
   fifo_reg_1_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n184, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_23_port);
   fifo_reg_1_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n182, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_22_port);
   fifo_reg_1_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n180, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_21_port);
   fifo_reg_1_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n178, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_20_port);
   fifo_reg_1_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n176, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_19_port);
   fifo_reg_1_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n174, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_18_port);
   fifo_reg_1_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n172, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_17_port);
   fifo_reg_1_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n170, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_16_port);
   fifo_reg_1_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n168, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_15_port);
   fifo_reg_1_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n166, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_14_port);
   fifo_reg_1_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n164, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_13_port);
   fifo_reg_1_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n162, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_12_port);
   fifo_reg_1_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n160, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_11_port);
   fifo_reg_1_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n158, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_1_10_port);
   fifo_reg_1_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n156, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_9_port);
   fifo_reg_1_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n154, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_8_port);
   fifo_reg_1_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n152, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_7_port);
   fifo_reg_1_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n150, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_6_port);
   fifo_reg_1_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n148, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_5_port);
   fifo_reg_1_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n146, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_1_4_port);
   fifo_reg_0_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n16, CLK => clk,
                           RESET => n45, SET => n1, QN => fifo_0_3_port);
   fifo_reg_0_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n14, CLK => clk,
                           RESET => n45, SET => n1, QN => fifo_0_2_port);
   fifo_reg_0_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n12, CLK => clk,
                           RESET => n45, SET => n1, QN => fifo_0_1_port);
   fifo_reg_0_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n10, CLK => clk,
                           RESET => n45, SET => n1, QN => fifo_0_0_port);
   fifo_reg_0_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n128, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_59_port);
   fifo_reg_0_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n126, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_58_port);
   fifo_reg_0_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n124, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_57_port);
   fifo_reg_0_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n122, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_56_port);
   fifo_reg_0_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n120, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_55_port);
   fifo_reg_0_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n118, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_54_port);
   fifo_reg_0_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n116, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_53_port);
   fifo_reg_0_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n114, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_52_port);
   fifo_reg_0_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n112, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_51_port);
   fifo_reg_0_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n110, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_50_port);
   fifo_reg_0_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n108, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_49_port);
   fifo_reg_0_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n106, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_48_port);
   fifo_reg_0_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n104, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_47_port);
   fifo_reg_0_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n102, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_46_port);
   fifo_reg_0_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n100, CLK => 
                           clk, RESET => n45, SET => n1, QN => fifo_0_45_port);
   fifo_reg_0_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n98, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_44_port);
   fifo_reg_0_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n96, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_43_port);
   fifo_reg_0_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n94, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_42_port);
   fifo_reg_0_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n92, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_41_port);
   fifo_reg_0_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n90, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_40_port);
   fifo_reg_0_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n88, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_39_port);
   fifo_reg_0_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n86, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_38_port);
   fifo_reg_0_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n84, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_37_port);
   fifo_reg_0_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n82, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_36_port);
   fifo_reg_0_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n80, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_35_port);
   fifo_reg_0_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n78, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_34_port);
   fifo_reg_0_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n76, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_33_port);
   fifo_reg_0_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n74, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_32_port);
   fifo_reg_0_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n72, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_31_port);
   fifo_reg_0_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n70, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_30_port);
   fifo_reg_0_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n68, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_29_port);
   fifo_reg_0_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n66, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_28_port);
   fifo_reg_0_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n64, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_27_port);
   fifo_reg_0_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n62, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_26_port);
   fifo_reg_0_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n60, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_25_port);
   fifo_reg_0_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n58, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_24_port);
   fifo_reg_0_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n56, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_23_port);
   fifo_reg_0_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n54, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_22_port);
   fifo_reg_0_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n52, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_21_port);
   fifo_reg_0_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n50, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_20_port);
   fifo_reg_0_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n48, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_19_port);
   fifo_reg_0_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n46, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_18_port);
   fifo_reg_0_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n44, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_17_port);
   fifo_reg_0_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n42, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_16_port);
   fifo_reg_0_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n40, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_15_port);
   fifo_reg_0_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n38, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_14_port);
   fifo_reg_0_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n36, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_13_port);
   fifo_reg_0_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n34, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_12_port);
   fifo_reg_0_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n32, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_11_port);
   fifo_reg_0_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n30, CLK => clk
                           , RESET => n45, SET => n1, QN => fifo_0_10_port);
   fifo_reg_0_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n28, CLK => clk,
                           RESET => n45, SET => n1, QN => fifo_0_9_port);
   fifo_reg_0_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n26, CLK => clk,
                           RESET => n45, SET => n1, QN => fifo_0_8_port);
   fifo_reg_0_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n24, CLK => clk,
                           RESET => n45, SET => n1, QN => fifo_0_7_port);
   fifo_reg_0_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n22, CLK => clk,
                           RESET => n45, SET => n1, QN => fifo_0_6_port);
   fifo_reg_0_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n20, CLK => clk,
                           RESET => n45, SET => n1, QN => fifo_0_5_port);
   fifo_reg_0_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n18, CLK => clk,
                           RESET => n45, SET => n1, QN => fifo_0_4_port);
   valid_data_reg : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n8, CLK => clk, 
                           RESET => n45, SET => n1, QN => valid_data_port);
   read_pointer_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n266, CLK 
                           => clk, RESET => n45, SET => n1, QN => 
                           read_pointer_0_port);
   U69 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U135 : INVx3_ASAP7_75t_R port map( A => rst, Y => n45);
   U138 : INVx1_ASAP7_75t_R port map( A => n29, Y => n17);
   U140 : INVx1_ASAP7_75t_R port map( A => n15, Y => n3);
   U141 : INVx1_ASAP7_75t_R port map( A => n31, Y => n43);
   U142 : HB1xp67_ASAP7_75t_R port map( A => n4, Y => n29);
   U207 : HB1xp67_ASAP7_75t_R port map( A => n6, Y => n15);
   U208 : HB1xp67_ASAP7_75t_R port map( A => n4, Y => n27);
   U209 : HB1xp67_ASAP7_75t_R port map( A => n4, Y => n25);
   U210 : HB1xp67_ASAP7_75t_R port map( A => n4, Y => n23);
   U211 : HB1xp67_ASAP7_75t_R port map( A => n4, Y => n21);
   U212 : HB1xp67_ASAP7_75t_R port map( A => n4, Y => n19);
   U213 : HB1xp67_ASAP7_75t_R port map( A => n6, Y => n13);
   U214 : HB1xp67_ASAP7_75t_R port map( A => n6, Y => n11);
   U215 : HB1xp67_ASAP7_75t_R port map( A => n6, Y => n9_port);
   U216 : HB1xp67_ASAP7_75t_R port map( A => n6, Y => n7_port);
   U217 : HB1xp67_ASAP7_75t_R port map( A => n6, Y => n5);
   U218 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n31);
   U219 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n33);
   U220 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n41);
   U221 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n39);
   U222 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n37);
   U223 : HB1xp67_ASAP7_75t_R port map( A => read_pointer_0_port, Y => n35);
   U224 : INVx1_ASAP7_75t_R port map( A => read_en, Y => n47);
   U225 : INVx1_ASAP7_75t_R port map( A => N7, Y => N9);
   U226 : INVx1_ASAP7_75t_R port map( A => write_en, Y => n49);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity arbiter_7_1_1_1_1_DXYU is

   port( clk, rst : in std_logic;  header : in std_logic_vector (129 downto 0);
         valid_data_vc_vec, incr_rx_vec : in std_logic_vector (12 downto 0);  
         crossbar_ctrl : out std_logic_vector (20 downto 0);  vc_transfer_vec, 
         vc_write_tx_vec : out std_logic_vector (12 downto 0));

end arbiter_7_1_1_1_1_DXYU;

architecture SYN_structural of arbiter_7_1_1_1_1_DXYU is

   component switch_allocator_7_DXYU
      port( clk, rst : in std_logic;  input_vc_in_use, output_vc_in_use : in 
            std_logic_vector (12 downto 0);  crossbar_ctrl_vec : in 
            std_logic_vector (38 downto 0);  vc_sel_enc_vec, valid_data_vc_vec,
            incr_rx_vec : in std_logic_vector (12 downto 0);  crossbar_ctrl : 
            out std_logic_vector (20 downto 0);  vc_transfer_vec, 
            vc_write_tx_vec : out std_logic_vector (12 downto 0));
   end component;
   
   component vc_allocator_7_1_1_1_1_DXYU
      port( clk, rst : in std_logic;  header : in std_logic_vector (129 downto 
            0);  enr_vc, valid_data_vc_vec : in std_logic_vector (12 downto 0);
            input_vc_in_use : out std_logic_vector (12 downto 0);  
            crossbar_ctrl_vec : out std_logic_vector (38 downto 0);  
            vc_sel_enc_vec, output_vc_in_use : out std_logic_vector (12 downto 
            0));
   end component;
   
   signal vc_transfer_vec_12_port, vc_transfer_vec_11_port, 
      vc_transfer_vec_10_port, vc_transfer_vec_9_port, vc_transfer_vec_8_port, 
      vc_transfer_vec_7_port, vc_transfer_vec_6_port, vc_transfer_vec_5_port, 
      vc_transfer_vec_4_port, vc_transfer_vec_3_port, vc_transfer_vec_2_port, 
      vc_transfer_vec_1_port, vc_transfer_vec_0_port, input_vc_in_use_12_port, 
      input_vc_in_use_11_port, input_vc_in_use_10_port, input_vc_in_use_9_port,
      input_vc_in_use_8_port, input_vc_in_use_7_port, input_vc_in_use_6_port, 
      input_vc_in_use_5_port, input_vc_in_use_4_port, input_vc_in_use_3_port, 
      input_vc_in_use_2_port, input_vc_in_use_1_port, input_vc_in_use_0_port, 
      crossbar_ctrl_vec_38_port, crossbar_ctrl_vec_37_port, 
      crossbar_ctrl_vec_36_port, crossbar_ctrl_vec_35_port, 
      crossbar_ctrl_vec_34_port, crossbar_ctrl_vec_33_port, 
      crossbar_ctrl_vec_32_port, crossbar_ctrl_vec_31_port, 
      crossbar_ctrl_vec_30_port, crossbar_ctrl_vec_29_port, 
      crossbar_ctrl_vec_28_port, crossbar_ctrl_vec_27_port, 
      crossbar_ctrl_vec_26_port, crossbar_ctrl_vec_25_port, 
      crossbar_ctrl_vec_24_port, crossbar_ctrl_vec_23_port, 
      crossbar_ctrl_vec_22_port, crossbar_ctrl_vec_21_port, 
      crossbar_ctrl_vec_20_port, crossbar_ctrl_vec_19_port, 
      crossbar_ctrl_vec_18_port, crossbar_ctrl_vec_17_port, 
      crossbar_ctrl_vec_16_port, crossbar_ctrl_vec_15_port, 
      crossbar_ctrl_vec_14_port, crossbar_ctrl_vec_13_port, 
      crossbar_ctrl_vec_12_port, crossbar_ctrl_vec_11_port, 
      crossbar_ctrl_vec_10_port, crossbar_ctrl_vec_9_port, 
      crossbar_ctrl_vec_8_port, crossbar_ctrl_vec_7_port, 
      crossbar_ctrl_vec_6_port, crossbar_ctrl_vec_5_port, 
      crossbar_ctrl_vec_4_port, crossbar_ctrl_vec_3_port, 
      crossbar_ctrl_vec_2_port, crossbar_ctrl_vec_1_port, 
      crossbar_ctrl_vec_0_port, vc_sel_enc_vec_12_0_port, 
      vc_sel_enc_vec_11_0_port, vc_sel_enc_vec_10_0_port, 
      vc_sel_enc_vec_9_0_port, vc_sel_enc_vec_8_0_port, vc_sel_enc_vec_7_0_port
      , vc_sel_enc_vec_6_0_port, vc_sel_enc_vec_5_0_port, 
      vc_sel_enc_vec_4_0_port, vc_sel_enc_vec_3_0_port, vc_sel_enc_vec_2_0_port
      , vc_sel_enc_vec_1_0_port, vc_sel_enc_vec_0_0_port, 
      output_vc_in_use_12_port, output_vc_in_use_11_port, 
      output_vc_in_use_10_port, output_vc_in_use_9_port, 
      output_vc_in_use_8_port, output_vc_in_use_7_port, output_vc_in_use_6_port
      , output_vc_in_use_5_port, output_vc_in_use_4_port, 
      output_vc_in_use_3_port, output_vc_in_use_2_port, output_vc_in_use_1_port
      , output_vc_in_use_0_port : std_logic;

begin
   vc_transfer_vec <= ( vc_transfer_vec_12_port, vc_transfer_vec_11_port, 
      vc_transfer_vec_10_port, vc_transfer_vec_9_port, vc_transfer_vec_8_port, 
      vc_transfer_vec_7_port, vc_transfer_vec_6_port, vc_transfer_vec_5_port, 
      vc_transfer_vec_4_port, vc_transfer_vec_3_port, vc_transfer_vec_2_port, 
      vc_transfer_vec_1_port, vc_transfer_vec_0_port );
   
   vc_allocator_1 : vc_allocator_7_1_1_1_1_DXYU port map( clk => clk, rst => 
                           rst, header(129) => header(129), header(128) => 
                           header(128), header(127) => header(127), header(126)
                           => header(126), header(125) => header(125), 
                           header(124) => header(124), header(123) => 
                           header(123), header(122) => header(122), header(121)
                           => header(121), header(120) => header(120), 
                           header(119) => header(119), header(118) => 
                           header(118), header(117) => header(117), header(116)
                           => header(116), header(115) => header(115), 
                           header(114) => header(114), header(113) => 
                           header(113), header(112) => header(112), header(111)
                           => header(111), header(110) => header(110), 
                           header(109) => header(109), header(108) => 
                           header(108), header(107) => header(107), header(106)
                           => header(106), header(105) => header(105), 
                           header(104) => header(104), header(103) => 
                           header(103), header(102) => header(102), header(101)
                           => header(101), header(100) => header(100), 
                           header(99) => header(99), header(98) => header(98), 
                           header(97) => header(97), header(96) => header(96), 
                           header(95) => header(95), header(94) => header(94), 
                           header(93) => header(93), header(92) => header(92), 
                           header(91) => header(91), header(90) => header(90), 
                           header(89) => header(89), header(88) => header(88), 
                           header(87) => header(87), header(86) => header(86), 
                           header(85) => header(85), header(84) => header(84), 
                           header(83) => header(83), header(82) => header(82), 
                           header(81) => header(81), header(80) => header(80), 
                           header(79) => header(79), header(78) => header(78), 
                           header(77) => header(77), header(76) => header(76), 
                           header(75) => header(75), header(74) => header(74), 
                           header(73) => header(73), header(72) => header(72), 
                           header(71) => header(71), header(70) => header(70), 
                           header(69) => header(69), header(68) => header(68), 
                           header(67) => header(67), header(66) => header(66), 
                           header(65) => header(65), header(64) => header(64), 
                           header(63) => header(63), header(62) => header(62), 
                           header(61) => header(61), header(60) => header(60), 
                           header(59) => header(59), header(58) => header(58), 
                           header(57) => header(57), header(56) => header(56), 
                           header(55) => header(55), header(54) => header(54), 
                           header(53) => header(53), header(52) => header(52), 
                           header(51) => header(51), header(50) => header(50), 
                           header(49) => header(49), header(48) => header(48), 
                           header(47) => header(47), header(46) => header(46), 
                           header(45) => header(45), header(44) => header(44), 
                           header(43) => header(43), header(42) => header(42), 
                           header(41) => header(41), header(40) => header(40), 
                           header(39) => header(39), header(38) => header(38), 
                           header(37) => header(37), header(36) => header(36), 
                           header(35) => header(35), header(34) => header(34), 
                           header(33) => header(33), header(32) => header(32), 
                           header(31) => header(31), header(30) => header(30), 
                           header(29) => header(29), header(28) => header(28), 
                           header(27) => header(27), header(26) => header(26), 
                           header(25) => header(25), header(24) => header(24), 
                           header(23) => header(23), header(22) => header(22), 
                           header(21) => header(21), header(20) => header(20), 
                           header(19) => header(19), header(18) => header(18), 
                           header(17) => header(17), header(16) => header(16), 
                           header(15) => header(15), header(14) => header(14), 
                           header(13) => header(13), header(12) => header(12), 
                           header(11) => header(11), header(10) => header(10), 
                           header(9) => header(9), header(8) => header(8), 
                           header(7) => header(7), header(6) => header(6), 
                           header(5) => header(5), header(4) => header(4), 
                           header(3) => header(3), header(2) => header(2), 
                           header(1) => header(1), header(0) => header(0), 
                           enr_vc(12) => vc_transfer_vec_12_port, enr_vc(11) =>
                           vc_transfer_vec_11_port, enr_vc(10) => 
                           vc_transfer_vec_10_port, enr_vc(9) => 
                           vc_transfer_vec_9_port, enr_vc(8) => 
                           vc_transfer_vec_8_port, enr_vc(7) => 
                           vc_transfer_vec_7_port, enr_vc(6) => 
                           vc_transfer_vec_6_port, enr_vc(5) => 
                           vc_transfer_vec_5_port, enr_vc(4) => 
                           vc_transfer_vec_4_port, enr_vc(3) => 
                           vc_transfer_vec_3_port, enr_vc(2) => 
                           vc_transfer_vec_2_port, enr_vc(1) => 
                           vc_transfer_vec_1_port, enr_vc(0) => 
                           vc_transfer_vec_0_port, valid_data_vc_vec(12) => 
                           valid_data_vc_vec(12), valid_data_vc_vec(11) => 
                           valid_data_vc_vec(11), valid_data_vc_vec(10) => 
                           valid_data_vc_vec(10), valid_data_vc_vec(9) => 
                           valid_data_vc_vec(9), valid_data_vc_vec(8) => 
                           valid_data_vc_vec(8), valid_data_vc_vec(7) => 
                           valid_data_vc_vec(7), valid_data_vc_vec(6) => 
                           valid_data_vc_vec(6), valid_data_vc_vec(5) => 
                           valid_data_vc_vec(5), valid_data_vc_vec(4) => 
                           valid_data_vc_vec(4), valid_data_vc_vec(3) => 
                           valid_data_vc_vec(3), valid_data_vc_vec(2) => 
                           valid_data_vc_vec(2), valid_data_vc_vec(1) => 
                           valid_data_vc_vec(1), valid_data_vc_vec(0) => 
                           valid_data_vc_vec(0), input_vc_in_use(12) => 
                           input_vc_in_use_12_port, input_vc_in_use(11) => 
                           input_vc_in_use_11_port, input_vc_in_use(10) => 
                           input_vc_in_use_10_port, input_vc_in_use(9) => 
                           input_vc_in_use_9_port, input_vc_in_use(8) => 
                           input_vc_in_use_8_port, input_vc_in_use(7) => 
                           input_vc_in_use_7_port, input_vc_in_use(6) => 
                           input_vc_in_use_6_port, input_vc_in_use(5) => 
                           input_vc_in_use_5_port, input_vc_in_use(4) => 
                           input_vc_in_use_4_port, input_vc_in_use(3) => 
                           input_vc_in_use_3_port, input_vc_in_use(2) => 
                           input_vc_in_use_2_port, input_vc_in_use(1) => 
                           input_vc_in_use_1_port, input_vc_in_use(0) => 
                           input_vc_in_use_0_port, crossbar_ctrl_vec(38) => 
                           crossbar_ctrl_vec_38_port, crossbar_ctrl_vec(37) => 
                           crossbar_ctrl_vec_37_port, crossbar_ctrl_vec(36) => 
                           crossbar_ctrl_vec_36_port, crossbar_ctrl_vec(35) => 
                           crossbar_ctrl_vec_35_port, crossbar_ctrl_vec(34) => 
                           crossbar_ctrl_vec_34_port, crossbar_ctrl_vec(33) => 
                           crossbar_ctrl_vec_33_port, crossbar_ctrl_vec(32) => 
                           crossbar_ctrl_vec_32_port, crossbar_ctrl_vec(31) => 
                           crossbar_ctrl_vec_31_port, crossbar_ctrl_vec(30) => 
                           crossbar_ctrl_vec_30_port, crossbar_ctrl_vec(29) => 
                           crossbar_ctrl_vec_29_port, crossbar_ctrl_vec(28) => 
                           crossbar_ctrl_vec_28_port, crossbar_ctrl_vec(27) => 
                           crossbar_ctrl_vec_27_port, crossbar_ctrl_vec(26) => 
                           crossbar_ctrl_vec_26_port, crossbar_ctrl_vec(25) => 
                           crossbar_ctrl_vec_25_port, crossbar_ctrl_vec(24) => 
                           crossbar_ctrl_vec_24_port, crossbar_ctrl_vec(23) => 
                           crossbar_ctrl_vec_23_port, crossbar_ctrl_vec(22) => 
                           crossbar_ctrl_vec_22_port, crossbar_ctrl_vec(21) => 
                           crossbar_ctrl_vec_21_port, crossbar_ctrl_vec(20) => 
                           crossbar_ctrl_vec_20_port, crossbar_ctrl_vec(19) => 
                           crossbar_ctrl_vec_19_port, crossbar_ctrl_vec(18) => 
                           crossbar_ctrl_vec_18_port, crossbar_ctrl_vec(17) => 
                           crossbar_ctrl_vec_17_port, crossbar_ctrl_vec(16) => 
                           crossbar_ctrl_vec_16_port, crossbar_ctrl_vec(15) => 
                           crossbar_ctrl_vec_15_port, crossbar_ctrl_vec(14) => 
                           crossbar_ctrl_vec_14_port, crossbar_ctrl_vec(13) => 
                           crossbar_ctrl_vec_13_port, crossbar_ctrl_vec(12) => 
                           crossbar_ctrl_vec_12_port, crossbar_ctrl_vec(11) => 
                           crossbar_ctrl_vec_11_port, crossbar_ctrl_vec(10) => 
                           crossbar_ctrl_vec_10_port, crossbar_ctrl_vec(9) => 
                           crossbar_ctrl_vec_9_port, crossbar_ctrl_vec(8) => 
                           crossbar_ctrl_vec_8_port, crossbar_ctrl_vec(7) => 
                           crossbar_ctrl_vec_7_port, crossbar_ctrl_vec(6) => 
                           crossbar_ctrl_vec_6_port, crossbar_ctrl_vec(5) => 
                           crossbar_ctrl_vec_5_port, crossbar_ctrl_vec(4) => 
                           crossbar_ctrl_vec_4_port, crossbar_ctrl_vec(3) => 
                           crossbar_ctrl_vec_3_port, crossbar_ctrl_vec(2) => 
                           crossbar_ctrl_vec_2_port, crossbar_ctrl_vec(1) => 
                           crossbar_ctrl_vec_1_port, crossbar_ctrl_vec(0) => 
                           crossbar_ctrl_vec_0_port, vc_sel_enc_vec(12) => 
                           vc_sel_enc_vec_12_0_port, vc_sel_enc_vec(11) => 
                           vc_sel_enc_vec_11_0_port, vc_sel_enc_vec(10) => 
                           vc_sel_enc_vec_10_0_port, vc_sel_enc_vec(9) => 
                           vc_sel_enc_vec_9_0_port, vc_sel_enc_vec(8) => 
                           vc_sel_enc_vec_8_0_port, vc_sel_enc_vec(7) => 
                           vc_sel_enc_vec_7_0_port, vc_sel_enc_vec(6) => 
                           vc_sel_enc_vec_6_0_port, vc_sel_enc_vec(5) => 
                           vc_sel_enc_vec_5_0_port, vc_sel_enc_vec(4) => 
                           vc_sel_enc_vec_4_0_port, vc_sel_enc_vec(3) => 
                           vc_sel_enc_vec_3_0_port, vc_sel_enc_vec(2) => 
                           vc_sel_enc_vec_2_0_port, vc_sel_enc_vec(1) => 
                           vc_sel_enc_vec_1_0_port, vc_sel_enc_vec(0) => 
                           vc_sel_enc_vec_0_0_port, output_vc_in_use(12) => 
                           output_vc_in_use_12_port, output_vc_in_use(11) => 
                           output_vc_in_use_11_port, output_vc_in_use(10) => 
                           output_vc_in_use_10_port, output_vc_in_use(9) => 
                           output_vc_in_use_9_port, output_vc_in_use(8) => 
                           output_vc_in_use_8_port, output_vc_in_use(7) => 
                           output_vc_in_use_7_port, output_vc_in_use(6) => 
                           output_vc_in_use_6_port, output_vc_in_use(5) => 
                           output_vc_in_use_5_port, output_vc_in_use(4) => 
                           output_vc_in_use_4_port, output_vc_in_use(3) => 
                           output_vc_in_use_3_port, output_vc_in_use(2) => 
                           output_vc_in_use_2_port, output_vc_in_use(1) => 
                           output_vc_in_use_1_port, output_vc_in_use(0) => 
                           output_vc_in_use_0_port);
   switch_allocator_1 : switch_allocator_7_DXYU port map( clk => clk, rst => 
                           rst, input_vc_in_use(12) => input_vc_in_use_12_port,
                           input_vc_in_use(11) => input_vc_in_use_11_port, 
                           input_vc_in_use(10) => input_vc_in_use_10_port, 
                           input_vc_in_use(9) => input_vc_in_use_9_port, 
                           input_vc_in_use(8) => input_vc_in_use_8_port, 
                           input_vc_in_use(7) => input_vc_in_use_7_port, 
                           input_vc_in_use(6) => input_vc_in_use_6_port, 
                           input_vc_in_use(5) => input_vc_in_use_5_port, 
                           input_vc_in_use(4) => input_vc_in_use_4_port, 
                           input_vc_in_use(3) => input_vc_in_use_3_port, 
                           input_vc_in_use(2) => input_vc_in_use_2_port, 
                           input_vc_in_use(1) => input_vc_in_use_1_port, 
                           input_vc_in_use(0) => input_vc_in_use_0_port, 
                           output_vc_in_use(12) => output_vc_in_use_12_port, 
                           output_vc_in_use(11) => output_vc_in_use_11_port, 
                           output_vc_in_use(10) => output_vc_in_use_10_port, 
                           output_vc_in_use(9) => output_vc_in_use_9_port, 
                           output_vc_in_use(8) => output_vc_in_use_8_port, 
                           output_vc_in_use(7) => output_vc_in_use_7_port, 
                           output_vc_in_use(6) => output_vc_in_use_6_port, 
                           output_vc_in_use(5) => output_vc_in_use_5_port, 
                           output_vc_in_use(4) => output_vc_in_use_4_port, 
                           output_vc_in_use(3) => output_vc_in_use_3_port, 
                           output_vc_in_use(2) => output_vc_in_use_2_port, 
                           output_vc_in_use(1) => output_vc_in_use_1_port, 
                           output_vc_in_use(0) => output_vc_in_use_0_port, 
                           crossbar_ctrl_vec(38) => crossbar_ctrl_vec_38_port, 
                           crossbar_ctrl_vec(37) => crossbar_ctrl_vec_37_port, 
                           crossbar_ctrl_vec(36) => crossbar_ctrl_vec_36_port, 
                           crossbar_ctrl_vec(35) => crossbar_ctrl_vec_35_port, 
                           crossbar_ctrl_vec(34) => crossbar_ctrl_vec_34_port, 
                           crossbar_ctrl_vec(33) => crossbar_ctrl_vec_33_port, 
                           crossbar_ctrl_vec(32) => crossbar_ctrl_vec_32_port, 
                           crossbar_ctrl_vec(31) => crossbar_ctrl_vec_31_port, 
                           crossbar_ctrl_vec(30) => crossbar_ctrl_vec_30_port, 
                           crossbar_ctrl_vec(29) => crossbar_ctrl_vec_29_port, 
                           crossbar_ctrl_vec(28) => crossbar_ctrl_vec_28_port, 
                           crossbar_ctrl_vec(27) => crossbar_ctrl_vec_27_port, 
                           crossbar_ctrl_vec(26) => crossbar_ctrl_vec_26_port, 
                           crossbar_ctrl_vec(25) => crossbar_ctrl_vec_25_port, 
                           crossbar_ctrl_vec(24) => crossbar_ctrl_vec_24_port, 
                           crossbar_ctrl_vec(23) => crossbar_ctrl_vec_23_port, 
                           crossbar_ctrl_vec(22) => crossbar_ctrl_vec_22_port, 
                           crossbar_ctrl_vec(21) => crossbar_ctrl_vec_21_port, 
                           crossbar_ctrl_vec(20) => crossbar_ctrl_vec_20_port, 
                           crossbar_ctrl_vec(19) => crossbar_ctrl_vec_19_port, 
                           crossbar_ctrl_vec(18) => crossbar_ctrl_vec_18_port, 
                           crossbar_ctrl_vec(17) => crossbar_ctrl_vec_17_port, 
                           crossbar_ctrl_vec(16) => crossbar_ctrl_vec_16_port, 
                           crossbar_ctrl_vec(15) => crossbar_ctrl_vec_15_port, 
                           crossbar_ctrl_vec(14) => crossbar_ctrl_vec_14_port, 
                           crossbar_ctrl_vec(13) => crossbar_ctrl_vec_13_port, 
                           crossbar_ctrl_vec(12) => crossbar_ctrl_vec_12_port, 
                           crossbar_ctrl_vec(11) => crossbar_ctrl_vec_11_port, 
                           crossbar_ctrl_vec(10) => crossbar_ctrl_vec_10_port, 
                           crossbar_ctrl_vec(9) => crossbar_ctrl_vec_9_port, 
                           crossbar_ctrl_vec(8) => crossbar_ctrl_vec_8_port, 
                           crossbar_ctrl_vec(7) => crossbar_ctrl_vec_7_port, 
                           crossbar_ctrl_vec(6) => crossbar_ctrl_vec_6_port, 
                           crossbar_ctrl_vec(5) => crossbar_ctrl_vec_5_port, 
                           crossbar_ctrl_vec(4) => crossbar_ctrl_vec_4_port, 
                           crossbar_ctrl_vec(3) => crossbar_ctrl_vec_3_port, 
                           crossbar_ctrl_vec(2) => crossbar_ctrl_vec_2_port, 
                           crossbar_ctrl_vec(1) => crossbar_ctrl_vec_1_port, 
                           crossbar_ctrl_vec(0) => crossbar_ctrl_vec_0_port, 
                           vc_sel_enc_vec(12) => vc_sel_enc_vec_12_0_port, 
                           vc_sel_enc_vec(11) => vc_sel_enc_vec_11_0_port, 
                           vc_sel_enc_vec(10) => vc_sel_enc_vec_10_0_port, 
                           vc_sel_enc_vec(9) => vc_sel_enc_vec_9_0_port, 
                           vc_sel_enc_vec(8) => vc_sel_enc_vec_8_0_port, 
                           vc_sel_enc_vec(7) => vc_sel_enc_vec_7_0_port, 
                           vc_sel_enc_vec(6) => vc_sel_enc_vec_6_0_port, 
                           vc_sel_enc_vec(5) => vc_sel_enc_vec_5_0_port, 
                           vc_sel_enc_vec(4) => vc_sel_enc_vec_4_0_port, 
                           vc_sel_enc_vec(3) => vc_sel_enc_vec_3_0_port, 
                           vc_sel_enc_vec(2) => vc_sel_enc_vec_2_0_port, 
                           vc_sel_enc_vec(1) => vc_sel_enc_vec_1_0_port, 
                           vc_sel_enc_vec(0) => vc_sel_enc_vec_0_0_port, 
                           valid_data_vc_vec(12) => valid_data_vc_vec(12), 
                           valid_data_vc_vec(11) => valid_data_vc_vec(11), 
                           valid_data_vc_vec(10) => valid_data_vc_vec(10), 
                           valid_data_vc_vec(9) => valid_data_vc_vec(9), 
                           valid_data_vc_vec(8) => valid_data_vc_vec(8), 
                           valid_data_vc_vec(7) => valid_data_vc_vec(7), 
                           valid_data_vc_vec(6) => valid_data_vc_vec(6), 
                           valid_data_vc_vec(5) => valid_data_vc_vec(5), 
                           valid_data_vc_vec(4) => valid_data_vc_vec(4), 
                           valid_data_vc_vec(3) => valid_data_vc_vec(3), 
                           valid_data_vc_vec(2) => valid_data_vc_vec(2), 
                           valid_data_vc_vec(1) => valid_data_vc_vec(1), 
                           valid_data_vc_vec(0) => valid_data_vc_vec(0), 
                           incr_rx_vec(12) => incr_rx_vec(12), incr_rx_vec(11) 
                           => incr_rx_vec(11), incr_rx_vec(10) => 
                           incr_rx_vec(10), incr_rx_vec(9) => incr_rx_vec(9), 
                           incr_rx_vec(8) => incr_rx_vec(8), incr_rx_vec(7) => 
                           incr_rx_vec(7), incr_rx_vec(6) => incr_rx_vec(6), 
                           incr_rx_vec(5) => incr_rx_vec(5), incr_rx_vec(4) => 
                           incr_rx_vec(4), incr_rx_vec(3) => incr_rx_vec(3), 
                           incr_rx_vec(2) => incr_rx_vec(2), incr_rx_vec(1) => 
                           incr_rx_vec(1), incr_rx_vec(0) => incr_rx_vec(0), 
                           crossbar_ctrl(20) => crossbar_ctrl(20), 
                           crossbar_ctrl(19) => crossbar_ctrl(19), 
                           crossbar_ctrl(18) => crossbar_ctrl(18), 
                           crossbar_ctrl(17) => crossbar_ctrl(17), 
                           crossbar_ctrl(16) => crossbar_ctrl(16), 
                           crossbar_ctrl(15) => crossbar_ctrl(15), 
                           crossbar_ctrl(14) => crossbar_ctrl(14), 
                           crossbar_ctrl(13) => crossbar_ctrl(13), 
                           crossbar_ctrl(12) => crossbar_ctrl(12), 
                           crossbar_ctrl(11) => crossbar_ctrl(11), 
                           crossbar_ctrl(10) => crossbar_ctrl(10), 
                           crossbar_ctrl(9) => crossbar_ctrl(9), 
                           crossbar_ctrl(8) => crossbar_ctrl(8), 
                           crossbar_ctrl(7) => crossbar_ctrl(7), 
                           crossbar_ctrl(6) => crossbar_ctrl(6), 
                           crossbar_ctrl(5) => crossbar_ctrl(5), 
                           crossbar_ctrl(4) => crossbar_ctrl(4), 
                           crossbar_ctrl(3) => crossbar_ctrl(3), 
                           crossbar_ctrl(2) => crossbar_ctrl(2), 
                           crossbar_ctrl(1) => crossbar_ctrl(1), 
                           crossbar_ctrl(0) => crossbar_ctrl(0), 
                           vc_transfer_vec(12) => vc_transfer_vec_12_port, 
                           vc_transfer_vec(11) => vc_transfer_vec_11_port, 
                           vc_transfer_vec(10) => vc_transfer_vec_10_port, 
                           vc_transfer_vec(9) => vc_transfer_vec_9_port, 
                           vc_transfer_vec(8) => vc_transfer_vec_8_port, 
                           vc_transfer_vec(7) => vc_transfer_vec_7_port, 
                           vc_transfer_vec(6) => vc_transfer_vec_6_port, 
                           vc_transfer_vec(5) => vc_transfer_vec_5_port, 
                           vc_transfer_vec(4) => vc_transfer_vec_4_port, 
                           vc_transfer_vec(3) => vc_transfer_vec_3_port, 
                           vc_transfer_vec(2) => vc_transfer_vec_2_port, 
                           vc_transfer_vec(1) => vc_transfer_vec_1_port, 
                           vc_transfer_vec(0) => vc_transfer_vec_0_port, 
                           vc_write_tx_vec(12) => vc_write_tx_vec(12), 
                           vc_write_tx_vec(11) => vc_write_tx_vec(11), 
                           vc_write_tx_vec(10) => vc_write_tx_vec(10), 
                           vc_write_tx_vec(9) => vc_write_tx_vec(9), 
                           vc_write_tx_vec(8) => vc_write_tx_vec(8), 
                           vc_write_tx_vec(7) => vc_write_tx_vec(7), 
                           vc_write_tx_vec(6) => vc_write_tx_vec(6), 
                           vc_write_tx_vec(5) => vc_write_tx_vec(5), 
                           vc_write_tx_vec(4) => vc_write_tx_vec(4), 
                           vc_write_tx_vec(3) => vc_write_tx_vec(3), 
                           vc_write_tx_vec(2) => vc_write_tx_vec(2), 
                           vc_write_tx_vec(1) => vc_write_tx_vec(1), 
                           vc_write_tx_vec(0) => vc_write_tx_vec(0));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity output_register_vc_num2_vc_num_out2_0 is

   port( clk, rst : in std_logic;  data_tx : in std_logic_vector (63 downto 0);
         vc_write_tx, incr_tx : in std_logic_vector (1 downto 0);  data_tx_pl :
         out std_logic_vector (63 downto 0);  vc_write_tx_pl, incr_tx_pl : out 
         std_logic_vector (1 downto 0));

end output_register_vc_num2_vc_num_out2_0;

architecture SYN_rtl of output_register_vc_num2_vc_num_out2_0 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx2_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal data_tx_pl_63_port, data_tx_pl_62_port, data_tx_pl_61_port, 
      data_tx_pl_60_port, data_tx_pl_59_port, data_tx_pl_58_port, 
      data_tx_pl_57_port, data_tx_pl_56_port, data_tx_pl_55_port, 
      data_tx_pl_54_port, data_tx_pl_53_port, data_tx_pl_52_port, 
      data_tx_pl_51_port, data_tx_pl_50_port, data_tx_pl_49_port, 
      data_tx_pl_48_port, data_tx_pl_47_port, data_tx_pl_46_port, 
      data_tx_pl_45_port, data_tx_pl_44_port, data_tx_pl_43_port, 
      data_tx_pl_42_port, data_tx_pl_41_port, data_tx_pl_40_port, 
      data_tx_pl_39_port, data_tx_pl_38_port, data_tx_pl_37_port, 
      data_tx_pl_36_port, data_tx_pl_35_port, data_tx_pl_34_port, 
      data_tx_pl_33_port, data_tx_pl_32_port, data_tx_pl_31_port, 
      data_tx_pl_30_port, data_tx_pl_29_port, data_tx_pl_28_port, 
      data_tx_pl_27_port, data_tx_pl_26_port, data_tx_pl_25_port, 
      data_tx_pl_24_port, data_tx_pl_23_port, data_tx_pl_22_port, 
      data_tx_pl_21_port, data_tx_pl_20_port, data_tx_pl_19_port, 
      data_tx_pl_18_port, data_tx_pl_17_port, data_tx_pl_16_port, 
      data_tx_pl_15_port, data_tx_pl_14_port, data_tx_pl_13_port, 
      data_tx_pl_12_port, data_tx_pl_11_port, data_tx_pl_10_port, 
      data_tx_pl_9_port, data_tx_pl_8_port, data_tx_pl_7_port, 
      data_tx_pl_6_port, data_tx_pl_5_port, data_tx_pl_4_port, 
      data_tx_pl_3_port, data_tx_pl_2_port, data_tx_pl_1_port, 
      data_tx_pl_0_port, n2, n7, n9, n11, n13, n15, n17, n19, n21, n23, n25, 
      n27, n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55
      , n57, n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, 
      n85, n87, n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, 
      n111, n113, n115, n117, n119, n121, n123, n125, n127, n129, n131, n133, 
      n1, n3, n4, n5, n6, n8, n10, n12, n14, n16, n18, n20, n22 : std_logic;

begin
   data_tx_pl <= ( data_tx_pl_63_port, data_tx_pl_62_port, data_tx_pl_61_port, 
      data_tx_pl_60_port, data_tx_pl_59_port, data_tx_pl_58_port, 
      data_tx_pl_57_port, data_tx_pl_56_port, data_tx_pl_55_port, 
      data_tx_pl_54_port, data_tx_pl_53_port, data_tx_pl_52_port, 
      data_tx_pl_51_port, data_tx_pl_50_port, data_tx_pl_49_port, 
      data_tx_pl_48_port, data_tx_pl_47_port, data_tx_pl_46_port, 
      data_tx_pl_45_port, data_tx_pl_44_port, data_tx_pl_43_port, 
      data_tx_pl_42_port, data_tx_pl_41_port, data_tx_pl_40_port, 
      data_tx_pl_39_port, data_tx_pl_38_port, data_tx_pl_37_port, 
      data_tx_pl_36_port, data_tx_pl_35_port, data_tx_pl_34_port, 
      data_tx_pl_33_port, data_tx_pl_32_port, data_tx_pl_31_port, 
      data_tx_pl_30_port, data_tx_pl_29_port, data_tx_pl_28_port, 
      data_tx_pl_27_port, data_tx_pl_26_port, data_tx_pl_25_port, 
      data_tx_pl_24_port, data_tx_pl_23_port, data_tx_pl_22_port, 
      data_tx_pl_21_port, data_tx_pl_20_port, data_tx_pl_19_port, 
      data_tx_pl_18_port, data_tx_pl_17_port, data_tx_pl_16_port, 
      data_tx_pl_15_port, data_tx_pl_14_port, data_tx_pl_13_port, 
      data_tx_pl_12_port, data_tx_pl_11_port, data_tx_pl_10_port, 
      data_tx_pl_9_port, data_tx_pl_8_port, data_tx_pl_7_port, 
      data_tx_pl_6_port, data_tx_pl_5_port, data_tx_pl_4_port, 
      data_tx_pl_3_port, data_tx_pl_2_port, data_tx_pl_1_port, 
      data_tx_pl_0_port );
   
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(0), A2 => n3, B1 => 
                           data_tx_pl_0_port, B2 => n12, Y => n7);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(1), A2 => n3, B1 => 
                           data_tx_pl_1_port, B2 => n12, Y => n9);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(2), A2 => n3, B1 => 
                           data_tx_pl_2_port, B2 => n12, Y => n11);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(3), A2 => n3, B1 => 
                           data_tx_pl_3_port, B2 => n12, Y => n13);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(4), A2 => n3, B1 => 
                           data_tx_pl_4_port, B2 => n10, Y => n15);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(5), A2 => n3, B1 => 
                           data_tx_pl_5_port, B2 => n10, Y => n17);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(6), A2 => n3, B1 => 
                           data_tx_pl_6_port, B2 => n10, Y => n19);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(7), A2 => n3, B1 => 
                           data_tx_pl_7_port, B2 => n10, Y => n21);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(8), A2 => n3, B1 => 
                           data_tx_pl_8_port, B2 => n10, Y => n23);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(9), A2 => n3, B1 => 
                           data_tx_pl_9_port, B2 => n10, Y => n25);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(10), A2 => n3, B1 => 
                           data_tx_pl_10_port, B2 => n10, Y => n27);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(11), A2 => n3, B1 => 
                           data_tx_pl_11_port, B2 => n10, Y => n29);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(12), A2 => n3, B1 => 
                           data_tx_pl_12_port, B2 => n10, Y => n31);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(13), A2 => n3, B1 => 
                           data_tx_pl_13_port, B2 => n10, Y => n33);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(14), A2 => n3, B1 => 
                           data_tx_pl_14_port, B2 => n10, Y => n35);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(15), A2 => n3, B1 => 
                           data_tx_pl_15_port, B2 => n10, Y => n37);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(16), A2 => n3, B1 => 
                           data_tx_pl_16_port, B2 => n8, Y => n39);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(17), A2 => n3, B1 => 
                           data_tx_pl_17_port, B2 => n8, Y => n41);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(18), A2 => n3, B1 => 
                           data_tx_pl_18_port, B2 => n8, Y => n43);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(19), A2 => n3, B1 => 
                           data_tx_pl_19_port, B2 => n8, Y => n45);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(20), A2 => n3, B1 => 
                           data_tx_pl_20_port, B2 => n8, Y => n47);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(21), A2 => n3, B1 => 
                           data_tx_pl_21_port, B2 => n8, Y => n49);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(22), A2 => n3, B1 => 
                           data_tx_pl_22_port, B2 => n8, Y => n51);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(23), A2 => n3, B1 => 
                           data_tx_pl_23_port, B2 => n8, Y => n53);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(24), A2 => n3, B1 => 
                           data_tx_pl_24_port, B2 => n8, Y => n55);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(25), A2 => n3, B1 => 
                           data_tx_pl_25_port, B2 => n8, Y => n57);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(26), A2 => n3, B1 => 
                           data_tx_pl_26_port, B2 => n8, Y => n59);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(27), A2 => n3, B1 => 
                           data_tx_pl_27_port, B2 => n8, Y => n61);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(28), A2 => n3, B1 => 
                           data_tx_pl_28_port, B2 => n6, Y => n63);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(29), A2 => n3, B1 => 
                           data_tx_pl_29_port, B2 => n6, Y => n65);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(30), A2 => n3, B1 => 
                           data_tx_pl_30_port, B2 => n6, Y => n67);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(31), A2 => n3, B1 => 
                           data_tx_pl_31_port, B2 => n6, Y => n69);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(32), A2 => n3, B1 => 
                           data_tx_pl_32_port, B2 => n6, Y => n71);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(33), A2 => n3, B1 => 
                           data_tx_pl_33_port, B2 => n6, Y => n73);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(34), A2 => n3, B1 => 
                           data_tx_pl_34_port, B2 => n6, Y => n75);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(35), A2 => n3, B1 => 
                           data_tx_pl_35_port, B2 => n6, Y => n77);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(36), A2 => n3, B1 => 
                           data_tx_pl_36_port, B2 => n6, Y => n79);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(37), A2 => n3, B1 => 
                           data_tx_pl_37_port, B2 => n6, Y => n81);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(38), A2 => n3, B1 => 
                           data_tx_pl_38_port, B2 => n6, Y => n83);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(39), A2 => n3, B1 => 
                           data_tx_pl_39_port, B2 => n6, Y => n85);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(40), A2 => n3, B1 => 
                           data_tx_pl_40_port, B2 => n5, Y => n87);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(41), A2 => n3, B1 => 
                           data_tx_pl_41_port, B2 => n5, Y => n89);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(42), A2 => n3, B1 => 
                           data_tx_pl_42_port, B2 => n5, Y => n91);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(43), A2 => n3, B1 => 
                           data_tx_pl_43_port, B2 => n5, Y => n93);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(44), A2 => n3, B1 => 
                           data_tx_pl_44_port, B2 => n5, Y => n95);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(45), A2 => n3, B1 => 
                           data_tx_pl_45_port, B2 => n5, Y => n97);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(46), A2 => n3, B1 => 
                           data_tx_pl_46_port, B2 => n5, Y => n99);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(47), A2 => n3, B1 => 
                           data_tx_pl_47_port, B2 => n5, Y => n101);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(48), A2 => n3, B1 => 
                           data_tx_pl_48_port, B2 => n5, Y => n103);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(49), A2 => n3, B1 => 
                           data_tx_pl_49_port, B2 => n5, Y => n105);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(50), A2 => n3, B1 => 
                           data_tx_pl_50_port, B2 => n5, Y => n107);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(51), A2 => n3, B1 => 
                           data_tx_pl_51_port, B2 => n5, Y => n109);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(52), A2 => n3, B1 => 
                           data_tx_pl_52_port, B2 => n4, Y => n111);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(53), A2 => n3, B1 => 
                           data_tx_pl_53_port, B2 => n4, Y => n113);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(54), A2 => n3, B1 => 
                           data_tx_pl_54_port, B2 => n4, Y => n115);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(55), A2 => n3, B1 => 
                           data_tx_pl_55_port, B2 => n4, Y => n117);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(56), A2 => n3, B1 => 
                           data_tx_pl_56_port, B2 => n4, Y => n119);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(57), A2 => n3, B1 => 
                           data_tx_pl_57_port, B2 => n4, Y => n121);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(58), A2 => n3, B1 => 
                           data_tx_pl_58_port, B2 => n4, Y => n123);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(59), A2 => n3, B1 => 
                           data_tx_pl_59_port, B2 => n4, Y => n125);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(60), A2 => n3, B1 => 
                           data_tx_pl_60_port, B2 => n4, Y => n127);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(61), A2 => n3, B1 => 
                           data_tx_pl_61_port, B2 => n4, Y => n129);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(62), A2 => n3, B1 => 
                           data_tx_pl_62_port, B2 => n4, Y => n131);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => data_tx(63), A2 => n3, B1 => 
                           data_tx_pl_63_port, B2 => n4, Y => n133);
   U68 : NAND2xp5_ASAP7_75t_R port map( A => n20, B => n22, Y => n2);
   vc_write_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n20, CLK
                           => clk, RESET => n16, SET => n1, QN => 
                           vc_write_tx_pl(1));
   vc_write_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n22, CLK
                           => clk, RESET => n16, SET => n1, QN => 
                           vc_write_tx_pl(0));
   incr_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n14, CLK => 
                           clk, RESET => n16, SET => n1, QN => incr_tx_pl(1));
   incr_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n18, CLK => 
                           clk, RESET => n16, SET => n1, QN => incr_tx_pl(0));
   data_tx_pl_reg_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_50_port);
   data_tx_pl_reg_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_49_port);
   data_tx_pl_reg_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_48_port);
   data_tx_pl_reg_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_47_port);
   data_tx_pl_reg_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_46_port);
   data_tx_pl_reg_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_45_port);
   data_tx_pl_reg_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_44_port);
   data_tx_pl_reg_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_43_port);
   data_tx_pl_reg_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_42_port);
   data_tx_pl_reg_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_41_port);
   data_tx_pl_reg_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_40_port);
   data_tx_pl_reg_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_39_port);
   data_tx_pl_reg_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_38_port);
   data_tx_pl_reg_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_37_port);
   data_tx_pl_reg_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_36_port);
   data_tx_pl_reg_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n77, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_35_port);
   data_tx_pl_reg_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n75, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_34_port);
   data_tx_pl_reg_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n73, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_33_port);
   data_tx_pl_reg_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n71, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_32_port);
   data_tx_pl_reg_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n69, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_31_port);
   data_tx_pl_reg_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n67, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_30_port);
   data_tx_pl_reg_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n31, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_12_port);
   data_tx_pl_reg_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n29, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_11_port);
   data_tx_pl_reg_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n27, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_10_port);
   data_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n7, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_0_port);
   data_tx_pl_reg_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n133, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_63_port);
   data_tx_pl_reg_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n131, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_62_port);
   data_tx_pl_reg_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n129, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_61_port);
   data_tx_pl_reg_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n127, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_60_port);
   data_tx_pl_reg_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n125, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_59_port);
   data_tx_pl_reg_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n123, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_58_port);
   data_tx_pl_reg_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n121, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_57_port);
   data_tx_pl_reg_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n119, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_56_port);
   data_tx_pl_reg_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n117, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_55_port);
   data_tx_pl_reg_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n115, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_54_port);
   data_tx_pl_reg_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_53_port);
   data_tx_pl_reg_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_52_port);
   data_tx_pl_reg_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_51_port);
   data_tx_pl_reg_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n65, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_29_port);
   data_tx_pl_reg_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n63, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_28_port);
   data_tx_pl_reg_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n61, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_27_port);
   data_tx_pl_reg_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n59, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_26_port);
   data_tx_pl_reg_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n57, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_25_port);
   data_tx_pl_reg_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n55, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_24_port);
   data_tx_pl_reg_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_23_port);
   data_tx_pl_reg_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_22_port);
   data_tx_pl_reg_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n49, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_21_port);
   data_tx_pl_reg_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n47, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_20_port);
   data_tx_pl_reg_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n45, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_19_port);
   data_tx_pl_reg_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n43, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_18_port);
   data_tx_pl_reg_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n41, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_17_port);
   data_tx_pl_reg_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n39, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_16_port);
   data_tx_pl_reg_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n37, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_15_port);
   data_tx_pl_reg_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n35, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_14_port);
   data_tx_pl_reg_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n33, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_13_port);
   data_tx_pl_reg_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n25, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_9_port);
   data_tx_pl_reg_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n23, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_8_port);
   data_tx_pl_reg_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n21, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_7_port);
   data_tx_pl_reg_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n19, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_6_port);
   data_tx_pl_reg_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n17, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_5_port);
   data_tx_pl_reg_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n15, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_4_port);
   data_tx_pl_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n13, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_3_port);
   data_tx_pl_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n11, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_2_port);
   data_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n9, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_1_port);
   U67 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U69 : INVx2_ASAP7_75t_R port map( A => rst, Y => n16);
   U70 : INVx1_ASAP7_75t_R port map( A => n12, Y => n3);
   U71 : HB1xp67_ASAP7_75t_R port map( A => n2, Y => n12);
   U72 : HB1xp67_ASAP7_75t_R port map( A => n2, Y => n10);
   U73 : HB1xp67_ASAP7_75t_R port map( A => n2, Y => n8);
   U74 : HB1xp67_ASAP7_75t_R port map( A => n2, Y => n6);
   U75 : HB1xp67_ASAP7_75t_R port map( A => n2, Y => n5);
   U76 : HB1xp67_ASAP7_75t_R port map( A => n2, Y => n4);
   U77 : INVx1_ASAP7_75t_R port map( A => incr_tx(1), Y => n14);
   U78 : INVx1_ASAP7_75t_R port map( A => incr_tx(0), Y => n18);
   U79 : INVx1_ASAP7_75t_R port map( A => vc_write_tx(1), Y => n20);
   U80 : INVx1_ASAP7_75t_R port map( A => vc_write_tx(0), Y => n22);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity output_register_vc_num1_vc_num_out1 is

   port( clk, rst : in std_logic;  data_tx : in std_logic_vector (63 downto 0);
         vc_write_tx, incr_tx : in std_logic;  data_tx_pl : out 
         std_logic_vector (63 downto 0);  vc_write_tx_pl, incr_tx_pl : out 
         std_logic);

end output_register_vc_num1_vc_num_out1;

architecture SYN_rtl of output_register_vc_num1_vc_num_out1 is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx2_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component TIELOx1_ASAP7_75t_R
      port( L : out std_logic);
   end component;
   
   component ASYNC_DFFHx1_ASAP7_75t_R
      port( D, CLK, RESET, SET : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal data_tx_pl_63_port, data_tx_pl_62_port, data_tx_pl_61_port, 
      data_tx_pl_60_port, data_tx_pl_59_port, data_tx_pl_58_port, 
      data_tx_pl_57_port, data_tx_pl_56_port, data_tx_pl_55_port, 
      data_tx_pl_54_port, data_tx_pl_53_port, data_tx_pl_52_port, 
      data_tx_pl_51_port, data_tx_pl_50_port, data_tx_pl_49_port, 
      data_tx_pl_48_port, data_tx_pl_47_port, data_tx_pl_46_port, 
      data_tx_pl_45_port, data_tx_pl_44_port, data_tx_pl_43_port, 
      data_tx_pl_42_port, data_tx_pl_41_port, data_tx_pl_40_port, 
      data_tx_pl_39_port, data_tx_pl_38_port, data_tx_pl_37_port, 
      data_tx_pl_36_port, data_tx_pl_35_port, data_tx_pl_34_port, 
      data_tx_pl_33_port, data_tx_pl_32_port, data_tx_pl_31_port, 
      data_tx_pl_30_port, data_tx_pl_29_port, data_tx_pl_28_port, 
      data_tx_pl_27_port, data_tx_pl_26_port, data_tx_pl_25_port, 
      data_tx_pl_24_port, data_tx_pl_23_port, data_tx_pl_22_port, 
      data_tx_pl_21_port, data_tx_pl_20_port, data_tx_pl_19_port, 
      data_tx_pl_18_port, data_tx_pl_17_port, data_tx_pl_16_port, 
      data_tx_pl_15_port, data_tx_pl_14_port, data_tx_pl_13_port, 
      data_tx_pl_12_port, data_tx_pl_11_port, data_tx_pl_10_port, 
      data_tx_pl_9_port, data_tx_pl_8_port, data_tx_pl_7_port, 
      data_tx_pl_6_port, data_tx_pl_5_port, data_tx_pl_4_port, 
      data_tx_pl_3_port, data_tx_pl_2_port, data_tx_pl_1_port, 
      data_tx_pl_0_port, n3, n5, n7, n9, n11, n13, n15, n17, n19, n21, n23, n25
      , n27, n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, 
      n55, n57, n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83
      , n85, n87, n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, 
      n111, n113, n115, n117, n119, n121, n123, n125, n127, n129, n1, n2, n4, 
      n6, n8, n10, n12, n14, n16, n18 : std_logic;

begin
   data_tx_pl <= ( data_tx_pl_63_port, data_tx_pl_62_port, data_tx_pl_61_port, 
      data_tx_pl_60_port, data_tx_pl_59_port, data_tx_pl_58_port, 
      data_tx_pl_57_port, data_tx_pl_56_port, data_tx_pl_55_port, 
      data_tx_pl_54_port, data_tx_pl_53_port, data_tx_pl_52_port, 
      data_tx_pl_51_port, data_tx_pl_50_port, data_tx_pl_49_port, 
      data_tx_pl_48_port, data_tx_pl_47_port, data_tx_pl_46_port, 
      data_tx_pl_45_port, data_tx_pl_44_port, data_tx_pl_43_port, 
      data_tx_pl_42_port, data_tx_pl_41_port, data_tx_pl_40_port, 
      data_tx_pl_39_port, data_tx_pl_38_port, data_tx_pl_37_port, 
      data_tx_pl_36_port, data_tx_pl_35_port, data_tx_pl_34_port, 
      data_tx_pl_33_port, data_tx_pl_32_port, data_tx_pl_31_port, 
      data_tx_pl_30_port, data_tx_pl_29_port, data_tx_pl_28_port, 
      data_tx_pl_27_port, data_tx_pl_26_port, data_tx_pl_25_port, 
      data_tx_pl_24_port, data_tx_pl_23_port, data_tx_pl_22_port, 
      data_tx_pl_21_port, data_tx_pl_20_port, data_tx_pl_19_port, 
      data_tx_pl_18_port, data_tx_pl_17_port, data_tx_pl_16_port, 
      data_tx_pl_15_port, data_tx_pl_14_port, data_tx_pl_13_port, 
      data_tx_pl_12_port, data_tx_pl_11_port, data_tx_pl_10_port, 
      data_tx_pl_9_port, data_tx_pl_8_port, data_tx_pl_7_port, 
      data_tx_pl_6_port, data_tx_pl_5_port, data_tx_pl_4_port, 
      data_tx_pl_3_port, data_tx_pl_2_port, data_tx_pl_1_port, 
      data_tx_pl_0_port );
   
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => n14, A2 => data_tx_pl_0_port, B1 
                           => data_tx(0), B2 => n2, Y => n3);
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => n14, A2 => data_tx_pl_1_port, B1 
                           => data_tx(1), B2 => n2, Y => n5);
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => n14, A2 => data_tx_pl_2_port, B1 
                           => data_tx(2), B2 => n2, Y => n7);
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => n14, A2 => data_tx_pl_3_port, B1 
                           => data_tx(3), B2 => n2, Y => n9);
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => n12, A2 => data_tx_pl_4_port, B1 
                           => data_tx(4), B2 => n2, Y => n11);
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => n12, A2 => data_tx_pl_5_port, B1 
                           => data_tx(5), B2 => n2, Y => n13);
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => n12, A2 => data_tx_pl_6_port, B1 
                           => data_tx(6), B2 => n2, Y => n15);
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => n12, A2 => data_tx_pl_7_port, B1 
                           => data_tx(7), B2 => n2, Y => n17);
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => n12, A2 => data_tx_pl_8_port, B1 
                           => data_tx(8), B2 => n2, Y => n19);
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => n12, A2 => data_tx_pl_9_port, B1 
                           => data_tx(9), B2 => n2, Y => n21);
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => n12, A2 => data_tx_pl_10_port, B1
                           => data_tx(10), B2 => n2, Y => n23);
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => n12, A2 => data_tx_pl_11_port, B1
                           => data_tx(11), B2 => n2, Y => n25);
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => n12, A2 => data_tx_pl_12_port, B1
                           => data_tx(12), B2 => n2, Y => n27);
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => n12, A2 => data_tx_pl_13_port, B1
                           => data_tx(13), B2 => n2, Y => n29);
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => n12, A2 => data_tx_pl_14_port, B1
                           => data_tx(14), B2 => n2, Y => n31);
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => n12, A2 => data_tx_pl_15_port, B1
                           => data_tx(15), B2 => n2, Y => n33);
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => n10, A2 => data_tx_pl_16_port, B1
                           => data_tx(16), B2 => n2, Y => n35);
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => n10, A2 => data_tx_pl_17_port, B1
                           => data_tx(17), B2 => n2, Y => n37);
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => n10, A2 => data_tx_pl_18_port, B1
                           => data_tx(18), B2 => n2, Y => n39);
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => n10, A2 => data_tx_pl_19_port, B1
                           => data_tx(19), B2 => n2, Y => n41);
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => n10, A2 => data_tx_pl_20_port, B1
                           => data_tx(20), B2 => n2, Y => n43);
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => n10, A2 => data_tx_pl_21_port, B1
                           => data_tx(21), B2 => n2, Y => n45);
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => n10, A2 => data_tx_pl_22_port, B1
                           => data_tx(22), B2 => n2, Y => n47);
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => n10, A2 => data_tx_pl_23_port, B1
                           => data_tx(23), B2 => n2, Y => n49);
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => n10, A2 => data_tx_pl_24_port, B1
                           => data_tx(24), B2 => n2, Y => n51);
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => n10, A2 => data_tx_pl_25_port, B1
                           => data_tx(25), B2 => n2, Y => n53);
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => n10, A2 => data_tx_pl_26_port, B1
                           => data_tx(26), B2 => n2, Y => n55);
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => n10, A2 => data_tx_pl_27_port, B1
                           => data_tx(27), B2 => n2, Y => n57);
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => n8, A2 => data_tx_pl_28_port, B1 
                           => data_tx(28), B2 => n2, Y => n59);
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => n8, A2 => data_tx_pl_29_port, B1 
                           => data_tx(29), B2 => n2, Y => n61);
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => n8, A2 => data_tx_pl_30_port, B1 
                           => data_tx(30), B2 => n2, Y => n63);
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => n8, A2 => data_tx_pl_31_port, B1 
                           => data_tx(31), B2 => n2, Y => n65);
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => n8, A2 => data_tx_pl_32_port, B1 
                           => data_tx(32), B2 => n2, Y => n67);
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => n8, A2 => data_tx_pl_33_port, B1 
                           => data_tx(33), B2 => n2, Y => n69);
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => n8, A2 => data_tx_pl_34_port, B1 
                           => data_tx(34), B2 => n2, Y => n71);
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => n8, A2 => data_tx_pl_35_port, B1 
                           => data_tx(35), B2 => n2, Y => n73);
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => n8, A2 => data_tx_pl_36_port, B1 
                           => data_tx(36), B2 => n2, Y => n75);
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => n8, A2 => data_tx_pl_37_port, B1 
                           => data_tx(37), B2 => n2, Y => n77);
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => n8, A2 => data_tx_pl_38_port, B1 
                           => data_tx(38), B2 => n2, Y => n79);
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => n8, A2 => data_tx_pl_39_port, B1 
                           => data_tx(39), B2 => n2, Y => n81);
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => n6, A2 => data_tx_pl_40_port, B1 
                           => data_tx(40), B2 => n2, Y => n83);
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => n6, A2 => data_tx_pl_41_port, B1 
                           => data_tx(41), B2 => n2, Y => n85);
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => n6, A2 => data_tx_pl_42_port, B1 
                           => data_tx(42), B2 => n2, Y => n87);
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => n6, A2 => data_tx_pl_43_port, B1 
                           => data_tx(43), B2 => n2, Y => n89);
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => n6, A2 => data_tx_pl_44_port, B1 
                           => data_tx(44), B2 => n2, Y => n91);
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => n6, A2 => data_tx_pl_45_port, B1 
                           => data_tx(45), B2 => n2, Y => n93);
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => n6, A2 => data_tx_pl_46_port, B1 
                           => data_tx(46), B2 => n2, Y => n95);
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => n6, A2 => data_tx_pl_47_port, B1 
                           => data_tx(47), B2 => n2, Y => n97);
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => n6, A2 => data_tx_pl_48_port, B1 
                           => data_tx(48), B2 => n2, Y => n99);
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => n6, A2 => data_tx_pl_49_port, B1 
                           => data_tx(49), B2 => n2, Y => n101);
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => n6, A2 => data_tx_pl_50_port, B1 
                           => data_tx(50), B2 => n2, Y => n103);
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => n6, A2 => data_tx_pl_51_port, B1 
                           => data_tx(51), B2 => n2, Y => n105);
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => n4, A2 => data_tx_pl_52_port, B1 
                           => data_tx(52), B2 => n2, Y => n107);
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => n4, A2 => data_tx_pl_53_port, B1 
                           => data_tx(53), B2 => n2, Y => n109);
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => n4, A2 => data_tx_pl_54_port, B1 
                           => data_tx(54), B2 => n2, Y => n111);
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => n4, A2 => data_tx_pl_55_port, B1 
                           => data_tx(55), B2 => n2, Y => n113);
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => n4, A2 => data_tx_pl_56_port, B1 
                           => data_tx(56), B2 => n2, Y => n115);
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => n4, A2 => data_tx_pl_57_port, B1 
                           => data_tx(57), B2 => n2, Y => n117);
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => n4, A2 => data_tx_pl_58_port, B1 
                           => data_tx(58), B2 => n2, Y => n119);
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => n4, A2 => data_tx_pl_59_port, B1 
                           => data_tx(59), B2 => n2, Y => n121);
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => n4, A2 => data_tx_pl_60_port, B1 
                           => data_tx(60), B2 => n2, Y => n123);
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => n4, A2 => data_tx_pl_61_port, B1 
                           => data_tx(61), B2 => n2, Y => n125);
   U65 : OAI22xp5_ASAP7_75t_R port map( A1 => n4, A2 => data_tx_pl_62_port, B1 
                           => data_tx(62), B2 => n2, Y => n127);
   U66 : OAI22xp5_ASAP7_75t_R port map( A1 => n4, A2 => data_tx_pl_63_port, B1 
                           => data_tx(63), B2 => n2, Y => n129);
   vc_write_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n2, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           vc_write_tx_pl);
   incr_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n18, CLK => 
                           clk, RESET => n16, SET => n1, QN => incr_tx_pl);
   data_tx_pl_reg_50_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n103, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_50_port);
   data_tx_pl_reg_49_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n101, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_49_port);
   data_tx_pl_reg_48_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n99, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_48_port);
   data_tx_pl_reg_47_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n97, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_47_port);
   data_tx_pl_reg_46_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n95, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_46_port);
   data_tx_pl_reg_45_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n93, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_45_port);
   data_tx_pl_reg_44_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n91, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_44_port);
   data_tx_pl_reg_43_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n89, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_43_port);
   data_tx_pl_reg_42_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n87, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_42_port);
   data_tx_pl_reg_41_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n85, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_41_port);
   data_tx_pl_reg_40_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n83, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_40_port);
   data_tx_pl_reg_39_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n81, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_39_port);
   data_tx_pl_reg_38_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n79, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_38_port);
   data_tx_pl_reg_37_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n77, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_37_port);
   data_tx_pl_reg_36_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n75, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_36_port);
   data_tx_pl_reg_35_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n73, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_35_port);
   data_tx_pl_reg_34_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n71, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_34_port);
   data_tx_pl_reg_33_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n69, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_33_port);
   data_tx_pl_reg_32_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n67, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_32_port);
   data_tx_pl_reg_31_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n65, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_31_port);
   data_tx_pl_reg_30_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n63, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_30_port);
   data_tx_pl_reg_12_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n27, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_12_port);
   data_tx_pl_reg_11_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n25, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_11_port);
   data_tx_pl_reg_10_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n23, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_10_port);
   data_tx_pl_reg_0_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n3, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_0_port);
   data_tx_pl_reg_9_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n21, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_9_port);
   data_tx_pl_reg_8_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n19, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_8_port);
   data_tx_pl_reg_7_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n17, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_7_port);
   data_tx_pl_reg_6_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n15, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_6_port);
   data_tx_pl_reg_5_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n13, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_5_port);
   data_tx_pl_reg_63_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n129, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_63_port);
   data_tx_pl_reg_62_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n127, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_62_port);
   data_tx_pl_reg_61_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n125, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_61_port);
   data_tx_pl_reg_60_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n123, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_60_port);
   data_tx_pl_reg_59_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n121, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_59_port);
   data_tx_pl_reg_58_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n119, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_58_port);
   data_tx_pl_reg_57_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n117, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_57_port);
   data_tx_pl_reg_51_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n105, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_51_port);
   data_tx_pl_reg_29_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n61, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_29_port);
   data_tx_pl_reg_28_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n59, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_28_port);
   data_tx_pl_reg_27_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n57, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_27_port);
   data_tx_pl_reg_26_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n55, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_26_port);
   data_tx_pl_reg_25_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n53, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_25_port);
   data_tx_pl_reg_24_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n51, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_24_port);
   data_tx_pl_reg_23_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n49, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_23_port);
   data_tx_pl_reg_22_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n47, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_22_port);
   data_tx_pl_reg_21_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n45, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_21_port);
   data_tx_pl_reg_20_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n43, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_20_port);
   data_tx_pl_reg_19_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n41, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_19_port);
   data_tx_pl_reg_18_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n39, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_18_port);
   data_tx_pl_reg_17_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n37, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_17_port);
   data_tx_pl_reg_16_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n35, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_16_port);
   data_tx_pl_reg_15_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n33, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_15_port);
   data_tx_pl_reg_14_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n31, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_14_port);
   data_tx_pl_reg_13_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n29, CLK =>
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_13_port);
   data_tx_pl_reg_4_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n11, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_4_port);
   data_tx_pl_reg_3_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n9, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_3_port);
   data_tx_pl_reg_2_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n7, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_2_port);
   data_tx_pl_reg_1_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n5, CLK => 
                           clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_1_port);
   data_tx_pl_reg_56_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n115, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_56_port);
   data_tx_pl_reg_55_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n113, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_55_port);
   data_tx_pl_reg_54_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n111, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_54_port);
   data_tx_pl_reg_53_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n109, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_53_port);
   data_tx_pl_reg_52_inst : ASYNC_DFFHx1_ASAP7_75t_R port map( D => n107, CLK 
                           => clk, RESET => n16, SET => n1, QN => 
                           data_tx_pl_52_port);
   U67 : TIELOx1_ASAP7_75t_R port map( L => n1);
   U68 : INVx2_ASAP7_75t_R port map( A => rst, Y => n16);
   U69 : INVx1_ASAP7_75t_R port map( A => n14, Y => n2);
   U70 : HB1xp67_ASAP7_75t_R port map( A => vc_write_tx, Y => n14);
   U71 : HB1xp67_ASAP7_75t_R port map( A => vc_write_tx, Y => n12);
   U72 : HB1xp67_ASAP7_75t_R port map( A => vc_write_tx, Y => n10);
   U73 : HB1xp67_ASAP7_75t_R port map( A => vc_write_tx, Y => n8);
   U74 : HB1xp67_ASAP7_75t_R port map( A => vc_write_tx, Y => n6);
   U75 : HB1xp67_ASAP7_75t_R port map( A => vc_write_tx, Y => n4);
   U76 : INVx1_ASAP7_75t_R port map( A => incr_tx, Y => n18);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity crossbar_7_DXYU is

   port( crossbar_in : in std_logic_vector (447 downto 0);  crossbar_ctrl : in 
         std_logic_vector (20 downto 0);  crossbar_out : out std_logic_vector 
         (447 downto 0));

end crossbar_7_DXYU;

architecture SYN_rtl of crossbar_7_DXYU is

   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2xp33_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3xp33_ASAP7_75t_R
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI222xp33_ASAP7_75t_R
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI211xp5_ASAP7_75t_R
      port( A1, A2, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI221xp5_ASAP7_75t_R
      port( A1, A2, B1, B2, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI222xp33_ASAP7_75t_R
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2xp5_ASAP7_75t_R
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22xp5_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, 
      n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, 
      n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, 
      n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, 
      n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, 
      n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, 
      n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, 
      n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, 
      n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, 
      n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, 
      n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, 
      n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, 
      n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, 
      n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, 
      n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, 
      n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, 
      n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, 
      n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, 
      n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, 
      n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, 
      n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, 
      n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, 
      n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, 
      n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, 
      n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, 
      n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, 
      n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, 
      n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, 
      n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, 
      n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, 
      n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
      n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
      n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, 
      n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, 
      n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, 
      n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
      n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, 
      n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, 
      n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, 
      n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, 
      n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, 
      n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, 
      n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, 
      n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, 
      n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, 
      n394, n395, n396, n397, n398, n399, n400, n401, n402, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
      n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
      n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n973, n974, n975, n976 : std_logic;

begin
   
   U1 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n320, B1 => n166, B2 
                           => n976, Y => crossbar_out(393));
   U2 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n321, B1 => n166, B2 
                           => n975, Y => crossbar_out(392));
   U3 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n322, B1 => n166, B2 
                           => n974, Y => crossbar_out(391));
   U4 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n323, B1 => n166, B2 
                           => n973, Y => crossbar_out(390));
   U5 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n330, B1 => n166, B2 
                           => n972, Y => crossbar_out(447));
   U6 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n331, B1 => n166, B2 
                           => n971, Y => crossbar_out(446));
   U7 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n332, B1 => n166, B2 
                           => n970, Y => crossbar_out(445));
   U8 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n333, B1 => n166, B2 
                           => n969, Y => crossbar_out(444));
   U9 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n324, B1 => n166, B2 
                           => n968, Y => crossbar_out(389));
   U10 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n334, B1 => n166, B2 
                           => n967, Y => crossbar_out(443));
   U11 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n335, B1 => n166, B2 
                           => n966, Y => crossbar_out(442));
   U12 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n336, B1 => n166, B2 
                           => n965, Y => crossbar_out(441));
   U13 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n337, B1 => n167, B2 
                           => n964, Y => crossbar_out(440));
   U14 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n338, B1 => n167, B2 
                           => n963, Y => crossbar_out(439));
   U15 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n339, B1 => n167, B2 
                           => n962, Y => crossbar_out(438));
   U16 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n340, B1 => n167, B2 
                           => n961, Y => crossbar_out(437));
   U17 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n341, B1 => n167, B2 
                           => n960, Y => crossbar_out(436));
   U18 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n342, B1 => n167, B2 
                           => n959, Y => crossbar_out(435));
   U19 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n343, B1 => n167, B2 
                           => n958, Y => crossbar_out(434));
   U20 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n325, B1 => n167, B2 
                           => n957, Y => crossbar_out(388));
   U21 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n344, B1 => n167, B2 
                           => n956, Y => crossbar_out(433));
   U22 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n345, B1 => n167, B2 
                           => n955, Y => crossbar_out(432));
   U23 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n346, B1 => n167, B2 
                           => n954, Y => crossbar_out(431));
   U24 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n347, B1 => n167, B2 
                           => n953, Y => crossbar_out(430));
   U25 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n348, B1 => n168, B2 
                           => n952, Y => crossbar_out(429));
   U26 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n349, B1 => n168, B2 
                           => n951, Y => crossbar_out(428));
   U27 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n350, B1 => n168, B2 
                           => n950, Y => crossbar_out(427));
   U28 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n351, B1 => n168, B2 
                           => n949, Y => crossbar_out(426));
   U29 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n352, B1 => n168, B2 
                           => n948, Y => crossbar_out(425));
   U30 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n353, B1 => n168, B2 
                           => n947, Y => crossbar_out(424));
   U31 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n326, B1 => n168, B2 
                           => n946, Y => crossbar_out(387));
   U32 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n354, B1 => n168, B2 
                           => n945, Y => crossbar_out(423));
   U33 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n355, B1 => n168, B2 
                           => n944, Y => crossbar_out(422));
   U34 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n356, B1 => n168, B2 
                           => n943, Y => crossbar_out(421));
   U35 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n357, B1 => n168, B2 
                           => n942, Y => crossbar_out(420));
   U36 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n358, B1 => n168, B2 
                           => n941, Y => crossbar_out(419));
   U37 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n359, B1 => n169, B2 
                           => n940, Y => crossbar_out(418));
   U38 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n360, B1 => n169, B2 
                           => n939, Y => crossbar_out(417));
   U39 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n361, B1 => n169, B2 
                           => n938, Y => crossbar_out(416));
   U40 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n362, B1 => n169, B2 
                           => n937, Y => crossbar_out(415));
   U41 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n363, B1 => n169, B2 
                           => n936, Y => crossbar_out(414));
   U42 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n327, B1 => n169, B2 
                           => n935, Y => crossbar_out(386));
   U43 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n300, B1 => n169, B2 
                           => n934, Y => crossbar_out(413));
   U44 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n301, B1 => n169, B2 
                           => n933, Y => crossbar_out(412));
   U45 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n302, B1 => n169, B2 
                           => n932, Y => crossbar_out(411));
   U46 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n303, B1 => n169, B2 
                           => n931, Y => crossbar_out(410));
   U47 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n304, B1 => n169, B2 
                           => n930, Y => crossbar_out(409));
   U48 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n305, B1 => n169, B2 
                           => n929, Y => crossbar_out(408));
   U49 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n306, B1 => n170, B2 
                           => n928, Y => crossbar_out(407));
   U50 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n307, B1 => n170, B2 
                           => n927, Y => crossbar_out(406));
   U51 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n308, B1 => n170, B2 
                           => n926, Y => crossbar_out(405));
   U52 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n309, B1 => n170, B2 
                           => n925, Y => crossbar_out(404));
   U53 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n328, B1 => n170, B2 
                           => n924, Y => crossbar_out(385));
   U54 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n310, B1 => n170, B2 
                           => n923, Y => crossbar_out(403));
   U55 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n311, B1 => n170, B2 
                           => n922, Y => crossbar_out(402));
   U56 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n312, B1 => n170, B2 
                           => n921, Y => crossbar_out(401));
   U57 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n313, B1 => n170, B2 
                           => n920, Y => crossbar_out(400));
   U58 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n314, B1 => n170, B2 
                           => n919, Y => crossbar_out(399));
   U59 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n315, B1 => n170, B2 
                           => n918, Y => crossbar_out(398));
   U60 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n316, B1 => n170, B2 
                           => n917, Y => crossbar_out(397));
   U61 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n317, B1 => n171, B2 
                           => n916, Y => crossbar_out(396));
   U62 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n318, B1 => n171, B2 
                           => n915, Y => crossbar_out(395));
   U63 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n319, B1 => n171, B2 
                           => n914, Y => crossbar_out(394));
   U64 : OAI22xp5_ASAP7_75t_R port map( A1 => n165, A2 => n329, B1 => n171, B2 
                           => n913, Y => crossbar_out(384));
   U65 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(73), A2 => n138, B1 
                           => n132, B2 => crossbar_in(9), Y => n404);
   U66 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(72), A2 => n138, B1 
                           => n132, B2 => crossbar_in(8), Y => n411);
   U67 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(71), A2 => n138, B1 
                           => n132, B2 => crossbar_in(7), Y => n413);
   U68 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(70), A2 => n138, B1 
                           => n132, B2 => crossbar_in(6), Y => n415);
   U69 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(127), A2 => n138, B1 
                           => n132, B2 => crossbar_in(63), Y => n417);
   U70 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(126), A2 => n138, B1 
                           => n132, B2 => crossbar_in(62), Y => n419);
   U71 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(125), A2 => n138, B1 
                           => n132, B2 => crossbar_in(61), Y => n421);
   U72 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(124), A2 => n138, B1 
                           => n132, B2 => crossbar_in(60), Y => n423);
   U73 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(69), A2 => n138, B1 
                           => n132, B2 => crossbar_in(5), Y => n425);
   U74 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(123), A2 => n138, B1 
                           => n132, B2 => crossbar_in(59), Y => n427);
   U75 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(122), A2 => n138, B1 
                           => n132, B2 => crossbar_in(58), Y => n429);
   U76 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(121), A2 => n138, B1 
                           => n132, B2 => crossbar_in(57), Y => n431);
   U77 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(120), A2 => n139, B1 
                           => n133, B2 => crossbar_in(56), Y => n433);
   U78 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(119), A2 => n139, B1 
                           => n133, B2 => crossbar_in(55), Y => n435);
   U79 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(118), A2 => n139, B1 
                           => n133, B2 => crossbar_in(54), Y => n437);
   U80 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(117), A2 => n139, B1 
                           => n133, B2 => crossbar_in(53), Y => n439);
   U81 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(116), A2 => n139, B1 
                           => n133, B2 => crossbar_in(52), Y => n441);
   U82 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(115), A2 => n139, B1 
                           => n133, B2 => crossbar_in(51), Y => n443);
   U83 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(114), A2 => n139, B1 
                           => n133, B2 => crossbar_in(50), Y => n445);
   U84 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(68), A2 => n139, B1 
                           => n133, B2 => crossbar_in(4), Y => n447);
   U85 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(113), A2 => n139, B1 
                           => n133, B2 => crossbar_in(49), Y => n449);
   U86 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(112), A2 => n139, B1 
                           => n133, B2 => crossbar_in(48), Y => n451);
   U87 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(111), A2 => n139, B1 
                           => n133, B2 => crossbar_in(47), Y => n453);
   U88 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(110), A2 => n139, B1 
                           => n133, B2 => crossbar_in(46), Y => n455);
   U89 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(109), A2 => n140, B1 
                           => n134, B2 => crossbar_in(45), Y => n457);
   U90 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(108), A2 => n140, B1 
                           => n134, B2 => crossbar_in(44), Y => n459);
   U91 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(107), A2 => n140, B1 
                           => n134, B2 => crossbar_in(43), Y => n461);
   U92 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(106), A2 => n140, B1 
                           => n134, B2 => crossbar_in(42), Y => n463);
   U93 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(105), A2 => n140, B1 
                           => n134, B2 => crossbar_in(41), Y => n465);
   U94 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(104), A2 => n140, B1 
                           => n134, B2 => crossbar_in(40), Y => n467);
   U95 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(67), A2 => n140, B1 
                           => n134, B2 => crossbar_in(3), Y => n469);
   U96 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(103), A2 => n140, B1 
                           => n134, B2 => crossbar_in(39), Y => n471);
   U97 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(102), A2 => n140, B1 
                           => n134, B2 => crossbar_in(38), Y => n473);
   U98 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(101), A2 => n140, B1 
                           => n134, B2 => crossbar_in(37), Y => n475);
   U99 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(100), A2 => n140, B1 
                           => n134, B2 => crossbar_in(36), Y => n477);
   U100 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(99), A2 => n140, B1 
                           => n134, B2 => crossbar_in(35), Y => n479);
   U101 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(98), A2 => n141, B1 
                           => n135, B2 => crossbar_in(34), Y => n481);
   U102 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(97), A2 => n141, B1 
                           => n135, B2 => crossbar_in(33), Y => n483);
   U103 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(96), A2 => n141, B1 
                           => n135, B2 => crossbar_in(32), Y => n485);
   U104 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(95), A2 => n141, B1 
                           => n135, B2 => crossbar_in(31), Y => n487);
   U105 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(94), A2 => n141, B1 
                           => n135, B2 => crossbar_in(30), Y => n489);
   U106 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(66), A2 => n141, B1 
                           => n135, B2 => crossbar_in(2), Y => n491);
   U107 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(93), A2 => n141, B1 
                           => n135, B2 => crossbar_in(29), Y => n493);
   U108 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(92), A2 => n141, B1 
                           => n135, B2 => crossbar_in(28), Y => n495);
   U109 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(91), A2 => n141, B1 
                           => n135, B2 => crossbar_in(27), Y => n497);
   U110 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(90), A2 => n141, B1 
                           => n135, B2 => crossbar_in(26), Y => n499);
   U111 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(89), A2 => n141, B1 
                           => n135, B2 => crossbar_in(25), Y => n501);
   U112 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(88), A2 => n141, B1 
                           => n135, B2 => crossbar_in(24), Y => n503);
   U113 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(87), A2 => n142, B1 
                           => n136, B2 => crossbar_in(23), Y => n505);
   U114 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(86), A2 => n142, B1 
                           => n136, B2 => crossbar_in(22), Y => n507);
   U115 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(85), A2 => n142, B1 
                           => n136, B2 => crossbar_in(21), Y => n509);
   U116 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(84), A2 => n142, B1 
                           => n136, B2 => crossbar_in(20), Y => n511);
   U117 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(65), A2 => n142, B1 
                           => n136, B2 => crossbar_in(1), Y => n513);
   U118 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(83), A2 => n142, B1 
                           => n136, B2 => crossbar_in(19), Y => n515);
   U119 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(82), A2 => n142, B1 
                           => n136, B2 => crossbar_in(18), Y => n517);
   U120 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(81), A2 => n142, B1 
                           => n136, B2 => crossbar_in(17), Y => n519);
   U121 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(80), A2 => n142, B1 
                           => n136, B2 => crossbar_in(16), Y => n521);
   U122 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(79), A2 => n142, B1 
                           => n136, B2 => crossbar_in(15), Y => n523);
   U123 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(78), A2 => n142, B1 
                           => n136, B2 => crossbar_in(14), Y => n525);
   U124 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(77), A2 => n142, B1 
                           => n136, B2 => crossbar_in(13), Y => n527);
   U125 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(76), A2 => n143, B1 
                           => n137, B2 => crossbar_in(12), Y => n529);
   U126 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(75), A2 => n143, B1 
                           => n137, B2 => crossbar_in(11), Y => n531);
   U127 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(74), A2 => n143, B1 
                           => n137, B2 => crossbar_in(10), Y => n533);
   U131 : AOI22xp5_ASAP7_75t_R port map( A1 => crossbar_in(64), A2 => n143, B1 
                           => n137, B2 => crossbar_in(0), Y => n535);
   U134 : NAND2xp5_ASAP7_75t_R port map( A => n18, B => n12, Y => n537);
   U138 : NAND2xp5_ASAP7_75t_R port map( A => n901, B => n902, Y => n538);
   U142 : NAND2xp5_ASAP7_75t_R port map( A => n907, B => n906, Y => n606);
   U143 : AOI22xp5_ASAP7_75t_R port map( A1 => n49, A2 => crossbar_in(201), B1 
                           => n43, B2 => crossbar_in(137), Y => n675);
   U144 : AOI22xp5_ASAP7_75t_R port map( A1 => n49, A2 => crossbar_in(200), B1 
                           => n43, B2 => crossbar_in(136), Y => n682);
   U145 : AOI22xp5_ASAP7_75t_R port map( A1 => n49, A2 => crossbar_in(199), B1 
                           => n43, B2 => crossbar_in(135), Y => n684);
   U146 : AOI22xp5_ASAP7_75t_R port map( A1 => n49, A2 => crossbar_in(198), B1 
                           => n43, B2 => crossbar_in(134), Y => n686);
   U147 : AOI22xp5_ASAP7_75t_R port map( A1 => n49, A2 => crossbar_in(255), B1 
                           => n43, B2 => crossbar_in(191), Y => n688);
   U148 : AOI22xp5_ASAP7_75t_R port map( A1 => n49, A2 => crossbar_in(254), B1 
                           => n43, B2 => crossbar_in(190), Y => n690);
   U149 : AOI22xp5_ASAP7_75t_R port map( A1 => n49, A2 => crossbar_in(253), B1 
                           => n43, B2 => crossbar_in(189), Y => n692);
   U150 : AOI22xp5_ASAP7_75t_R port map( A1 => n49, A2 => crossbar_in(252), B1 
                           => n43, B2 => crossbar_in(188), Y => n694);
   U151 : AOI22xp5_ASAP7_75t_R port map( A1 => n49, A2 => crossbar_in(197), B1 
                           => n43, B2 => crossbar_in(133), Y => n696);
   U152 : AOI22xp5_ASAP7_75t_R port map( A1 => n49, A2 => crossbar_in(251), B1 
                           => n43, B2 => crossbar_in(187), Y => n698);
   U153 : AOI22xp5_ASAP7_75t_R port map( A1 => n49, A2 => crossbar_in(250), B1 
                           => n43, B2 => crossbar_in(186), Y => n700);
   U154 : AOI22xp5_ASAP7_75t_R port map( A1 => n49, A2 => crossbar_in(249), B1 
                           => n43, B2 => crossbar_in(185), Y => n702);
   U155 : AOI22xp5_ASAP7_75t_R port map( A1 => n50, A2 => crossbar_in(248), B1 
                           => n44, B2 => crossbar_in(184), Y => n704);
   U156 : AOI22xp5_ASAP7_75t_R port map( A1 => n50, A2 => crossbar_in(247), B1 
                           => n44, B2 => crossbar_in(183), Y => n706);
   U157 : AOI22xp5_ASAP7_75t_R port map( A1 => n50, A2 => crossbar_in(246), B1 
                           => n44, B2 => crossbar_in(182), Y => n708);
   U158 : AOI22xp5_ASAP7_75t_R port map( A1 => n50, A2 => crossbar_in(245), B1 
                           => n44, B2 => crossbar_in(181), Y => n710);
   U159 : AOI22xp5_ASAP7_75t_R port map( A1 => n50, A2 => crossbar_in(244), B1 
                           => n44, B2 => crossbar_in(180), Y => n712);
   U160 : AOI22xp5_ASAP7_75t_R port map( A1 => n50, A2 => crossbar_in(243), B1 
                           => n44, B2 => crossbar_in(179), Y => n714);
   U161 : AOI22xp5_ASAP7_75t_R port map( A1 => n50, A2 => crossbar_in(242), B1 
                           => n44, B2 => crossbar_in(178), Y => n716);
   U162 : AOI22xp5_ASAP7_75t_R port map( A1 => n50, A2 => crossbar_in(196), B1 
                           => n44, B2 => crossbar_in(132), Y => n718);
   U163 : AOI22xp5_ASAP7_75t_R port map( A1 => n50, A2 => crossbar_in(241), B1 
                           => n44, B2 => crossbar_in(177), Y => n720);
   U164 : AOI22xp5_ASAP7_75t_R port map( A1 => n50, A2 => crossbar_in(240), B1 
                           => n44, B2 => crossbar_in(176), Y => n722);
   U165 : AOI22xp5_ASAP7_75t_R port map( A1 => n50, A2 => crossbar_in(239), B1 
                           => n44, B2 => crossbar_in(175), Y => n724);
   U166 : AOI22xp5_ASAP7_75t_R port map( A1 => n50, A2 => crossbar_in(238), B1 
                           => n44, B2 => crossbar_in(174), Y => n726);
   U167 : AOI22xp5_ASAP7_75t_R port map( A1 => n51, A2 => crossbar_in(237), B1 
                           => n45, B2 => crossbar_in(173), Y => n728);
   U168 : AOI22xp5_ASAP7_75t_R port map( A1 => n51, A2 => crossbar_in(236), B1 
                           => n45, B2 => crossbar_in(172), Y => n730);
   U169 : AOI22xp5_ASAP7_75t_R port map( A1 => n51, A2 => crossbar_in(235), B1 
                           => n45, B2 => crossbar_in(171), Y => n732);
   U170 : AOI22xp5_ASAP7_75t_R port map( A1 => n51, A2 => crossbar_in(234), B1 
                           => n45, B2 => crossbar_in(170), Y => n734);
   U171 : AOI22xp5_ASAP7_75t_R port map( A1 => n51, A2 => crossbar_in(233), B1 
                           => n45, B2 => crossbar_in(169), Y => n736);
   U172 : AOI22xp5_ASAP7_75t_R port map( A1 => n51, A2 => crossbar_in(232), B1 
                           => n45, B2 => crossbar_in(168), Y => n738);
   U173 : AOI22xp5_ASAP7_75t_R port map( A1 => n51, A2 => crossbar_in(195), B1 
                           => n45, B2 => crossbar_in(131), Y => n740);
   U174 : AOI22xp5_ASAP7_75t_R port map( A1 => n51, A2 => crossbar_in(231), B1 
                           => n45, B2 => crossbar_in(167), Y => n742);
   U175 : AOI22xp5_ASAP7_75t_R port map( A1 => n51, A2 => crossbar_in(230), B1 
                           => n45, B2 => crossbar_in(166), Y => n744);
   U176 : AOI22xp5_ASAP7_75t_R port map( A1 => n51, A2 => crossbar_in(229), B1 
                           => n45, B2 => crossbar_in(165), Y => n746);
   U177 : AOI22xp5_ASAP7_75t_R port map( A1 => n51, A2 => crossbar_in(228), B1 
                           => n45, B2 => crossbar_in(164), Y => n748);
   U178 : AOI22xp5_ASAP7_75t_R port map( A1 => n51, A2 => crossbar_in(227), B1 
                           => n45, B2 => crossbar_in(163), Y => n750);
   U179 : AOI22xp5_ASAP7_75t_R port map( A1 => n52, A2 => crossbar_in(226), B1 
                           => n46, B2 => crossbar_in(162), Y => n752);
   U180 : AOI22xp5_ASAP7_75t_R port map( A1 => n52, A2 => crossbar_in(225), B1 
                           => n46, B2 => crossbar_in(161), Y => n754);
   U181 : AOI22xp5_ASAP7_75t_R port map( A1 => n52, A2 => crossbar_in(224), B1 
                           => n46, B2 => crossbar_in(160), Y => n756);
   U182 : AOI22xp5_ASAP7_75t_R port map( A1 => n52, A2 => crossbar_in(223), B1 
                           => n46, B2 => crossbar_in(159), Y => n758);
   U183 : AOI22xp5_ASAP7_75t_R port map( A1 => n52, A2 => crossbar_in(222), B1 
                           => n46, B2 => crossbar_in(158), Y => n760);
   U184 : AOI22xp5_ASAP7_75t_R port map( A1 => n52, A2 => crossbar_in(194), B1 
                           => n46, B2 => crossbar_in(130), Y => n762);
   U185 : AOI22xp5_ASAP7_75t_R port map( A1 => n52, A2 => crossbar_in(221), B1 
                           => n46, B2 => crossbar_in(157), Y => n764);
   U186 : AOI22xp5_ASAP7_75t_R port map( A1 => n52, A2 => crossbar_in(220), B1 
                           => n46, B2 => crossbar_in(156), Y => n766);
   U187 : AOI22xp5_ASAP7_75t_R port map( A1 => n52, A2 => crossbar_in(219), B1 
                           => n46, B2 => crossbar_in(155), Y => n768);
   U188 : AOI22xp5_ASAP7_75t_R port map( A1 => n52, A2 => crossbar_in(218), B1 
                           => n46, B2 => crossbar_in(154), Y => n770);
   U189 : AOI22xp5_ASAP7_75t_R port map( A1 => n52, A2 => crossbar_in(217), B1 
                           => n46, B2 => crossbar_in(153), Y => n772);
   U190 : AOI22xp5_ASAP7_75t_R port map( A1 => n52, A2 => crossbar_in(216), B1 
                           => n46, B2 => crossbar_in(152), Y => n774);
   U191 : AOI22xp5_ASAP7_75t_R port map( A1 => n53, A2 => crossbar_in(215), B1 
                           => n47, B2 => crossbar_in(151), Y => n776);
   U192 : AOI22xp5_ASAP7_75t_R port map( A1 => n53, A2 => crossbar_in(214), B1 
                           => n47, B2 => crossbar_in(150), Y => n778);
   U193 : AOI22xp5_ASAP7_75t_R port map( A1 => n53, A2 => crossbar_in(213), B1 
                           => n47, B2 => crossbar_in(149), Y => n780);
   U194 : AOI22xp5_ASAP7_75t_R port map( A1 => n53, A2 => crossbar_in(212), B1 
                           => n47, B2 => crossbar_in(148), Y => n782);
   U195 : AOI22xp5_ASAP7_75t_R port map( A1 => n53, A2 => crossbar_in(193), B1 
                           => n47, B2 => crossbar_in(129), Y => n784);
   U196 : AOI22xp5_ASAP7_75t_R port map( A1 => n53, A2 => crossbar_in(211), B1 
                           => n47, B2 => crossbar_in(147), Y => n786);
   U197 : AOI22xp5_ASAP7_75t_R port map( A1 => n53, A2 => crossbar_in(210), B1 
                           => n47, B2 => crossbar_in(146), Y => n788);
   U198 : AOI22xp5_ASAP7_75t_R port map( A1 => n53, A2 => crossbar_in(209), B1 
                           => n47, B2 => crossbar_in(145), Y => n790);
   U199 : AOI22xp5_ASAP7_75t_R port map( A1 => n53, A2 => crossbar_in(208), B1 
                           => n47, B2 => crossbar_in(144), Y => n792);
   U200 : AOI22xp5_ASAP7_75t_R port map( A1 => n53, A2 => crossbar_in(207), B1 
                           => n47, B2 => crossbar_in(143), Y => n794);
   U201 : AOI22xp5_ASAP7_75t_R port map( A1 => n53, A2 => crossbar_in(206), B1 
                           => n47, B2 => crossbar_in(142), Y => n796);
   U202 : AOI22xp5_ASAP7_75t_R port map( A1 => n53, A2 => crossbar_in(205), B1 
                           => n47, B2 => crossbar_in(141), Y => n798);
   U203 : AOI22xp5_ASAP7_75t_R port map( A1 => n54, A2 => crossbar_in(204), B1 
                           => n48, B2 => crossbar_in(140), Y => n800);
   U204 : AOI22xp5_ASAP7_75t_R port map( A1 => n54, A2 => crossbar_in(203), B1 
                           => n48, B2 => crossbar_in(139), Y => n802);
   U205 : AOI22xp5_ASAP7_75t_R port map( A1 => n54, A2 => crossbar_in(202), B1 
                           => n48, B2 => crossbar_in(138), Y => n804);
   U209 : AOI22xp5_ASAP7_75t_R port map( A1 => n54, A2 => crossbar_in(192), B1 
                           => n48, B2 => crossbar_in(128), Y => n806);
   U614 : OAI211xp5_ASAP7_75t_R port map( A1 => n163, A2 => n384, B => n404, C 
                           => n405, Y => crossbar_out(329));
   U615 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(137), A2 => n154, 
                           B1 => crossbar_in(265), B2 => n149, C1 => 
                           crossbar_in(201), C2 => n144, Y => n405);
   U616 : OAI211xp5_ASAP7_75t_R port map( A1 => n163, A2 => n385, B => n411, C 
                           => n412, Y => crossbar_out(328));
   U617 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(136), A2 => n154, 
                           B1 => crossbar_in(264), B2 => n149, C1 => 
                           crossbar_in(200), C2 => n144, Y => n412);
   U618 : OAI211xp5_ASAP7_75t_R port map( A1 => n163, A2 => n386, B => n413, C 
                           => n414, Y => crossbar_out(327));
   U619 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(135), A2 => n154, 
                           B1 => crossbar_in(263), B2 => n149, C1 => 
                           crossbar_in(199), C2 => n144, Y => n414);
   U620 : OAI211xp5_ASAP7_75t_R port map( A1 => n163, A2 => n387, B => n415, C 
                           => n416, Y => crossbar_out(326));
   U621 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(134), A2 => n154, 
                           B1 => crossbar_in(262), B2 => n149, C1 => 
                           crossbar_in(198), C2 => n144, Y => n416);
   U622 : OAI211xp5_ASAP7_75t_R port map( A1 => n163, A2 => n394, B => n417, C 
                           => n418, Y => crossbar_out(383));
   U623 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(191), A2 => n154, 
                           B1 => crossbar_in(319), B2 => n149, C1 => 
                           crossbar_in(255), C2 => n144, Y => n418);
   U624 : OAI211xp5_ASAP7_75t_R port map( A1 => n163, A2 => n395, B => n419, C 
                           => n420, Y => crossbar_out(382));
   U625 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(190), A2 => n154, 
                           B1 => crossbar_in(318), B2 => n149, C1 => 
                           crossbar_in(254), C2 => n144, Y => n420);
   U626 : OAI211xp5_ASAP7_75t_R port map( A1 => n163, A2 => n396, B => n421, C 
                           => n422, Y => crossbar_out(381));
   U627 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(189), A2 => n154, 
                           B1 => crossbar_in(317), B2 => n149, C1 => 
                           crossbar_in(253), C2 => n144, Y => n422);
   U628 : OAI211xp5_ASAP7_75t_R port map( A1 => n163, A2 => n397, B => n423, C 
                           => n424, Y => crossbar_out(380));
   U629 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(188), A2 => n154, 
                           B1 => crossbar_in(316), B2 => n149, C1 => 
                           crossbar_in(252), C2 => n144, Y => n424);
   U630 : OAI211xp5_ASAP7_75t_R port map( A1 => n163, A2 => n388, B => n425, C 
                           => n426, Y => crossbar_out(325));
   U631 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(133), A2 => n154, 
                           B1 => crossbar_in(261), B2 => n149, C1 => 
                           crossbar_in(197), C2 => n144, Y => n426);
   U632 : OAI211xp5_ASAP7_75t_R port map( A1 => n163, A2 => n398, B => n427, C 
                           => n428, Y => crossbar_out(379));
   U633 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(187), A2 => n154, 
                           B1 => crossbar_in(315), B2 => n149, C1 => 
                           crossbar_in(251), C2 => n144, Y => n428);
   U634 : OAI211xp5_ASAP7_75t_R port map( A1 => n163, A2 => n399, B => n429, C 
                           => n430, Y => crossbar_out(378));
   U635 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(186), A2 => n154, 
                           B1 => crossbar_in(314), B2 => n149, C1 => 
                           crossbar_in(250), C2 => n144, Y => n430);
   U636 : OAI211xp5_ASAP7_75t_R port map( A1 => n163, A2 => n400, B => n431, C 
                           => n432, Y => crossbar_out(377));
   U637 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(185), A2 => n154, 
                           B1 => crossbar_in(313), B2 => n149, C1 => 
                           crossbar_in(249), C2 => n144, Y => n432);
   U638 : OAI211xp5_ASAP7_75t_R port map( A1 => n162, A2 => n401, B => n433, C 
                           => n434, Y => crossbar_out(376));
   U639 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(184), A2 => n154, 
                           B1 => crossbar_in(312), B2 => n149, C1 => 
                           crossbar_in(248), C2 => n144, Y => n434);
   U640 : OAI211xp5_ASAP7_75t_R port map( A1 => n162, A2 => n402, B => n435, C 
                           => n436, Y => crossbar_out(375));
   U641 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(183), A2 => n155, 
                           B1 => crossbar_in(311), B2 => n150, C1 => 
                           crossbar_in(247), C2 => n145, Y => n436);
   U642 : OAI211xp5_ASAP7_75t_R port map( A1 => n162, A2 => n808, B => n437, C 
                           => n438, Y => crossbar_out(374));
   U643 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(182), A2 => n155, 
                           B1 => crossbar_in(310), B2 => n150, C1 => 
                           crossbar_in(246), C2 => n145, Y => n438);
   U644 : OAI211xp5_ASAP7_75t_R port map( A1 => n162, A2 => n809, B => n439, C 
                           => n440, Y => crossbar_out(373));
   U645 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(181), A2 => n155, 
                           B1 => crossbar_in(309), B2 => n150, C1 => 
                           crossbar_in(245), C2 => n145, Y => n440);
   U646 : OAI211xp5_ASAP7_75t_R port map( A1 => n162, A2 => n810, B => n441, C 
                           => n442, Y => crossbar_out(372));
   U647 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(180), A2 => n155, 
                           B1 => crossbar_in(308), B2 => n150, C1 => 
                           crossbar_in(244), C2 => n145, Y => n442);
   U648 : OAI211xp5_ASAP7_75t_R port map( A1 => n162, A2 => n811, B => n443, C 
                           => n444, Y => crossbar_out(371));
   U649 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(179), A2 => n155, 
                           B1 => crossbar_in(307), B2 => n150, C1 => 
                           crossbar_in(243), C2 => n145, Y => n444);
   U650 : OAI211xp5_ASAP7_75t_R port map( A1 => n162, A2 => n812, B => n445, C 
                           => n446, Y => crossbar_out(370));
   U651 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(178), A2 => n155, 
                           B1 => crossbar_in(306), B2 => n150, C1 => 
                           crossbar_in(242), C2 => n145, Y => n446);
   U652 : OAI211xp5_ASAP7_75t_R port map( A1 => n162, A2 => n389, B => n447, C 
                           => n448, Y => crossbar_out(324));
   U653 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(132), A2 => n155, 
                           B1 => crossbar_in(260), B2 => n150, C1 => 
                           crossbar_in(196), C2 => n145, Y => n448);
   U654 : OAI211xp5_ASAP7_75t_R port map( A1 => n162, A2 => n813, B => n449, C 
                           => n450, Y => crossbar_out(369));
   U655 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(177), A2 => n155, 
                           B1 => crossbar_in(305), B2 => n150, C1 => 
                           crossbar_in(241), C2 => n145, Y => n450);
   U656 : OAI211xp5_ASAP7_75t_R port map( A1 => n162, A2 => n814, B => n451, C 
                           => n452, Y => crossbar_out(368));
   U657 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(176), A2 => n155, 
                           B1 => crossbar_in(304), B2 => n150, C1 => 
                           crossbar_in(240), C2 => n145, Y => n452);
   U658 : OAI211xp5_ASAP7_75t_R port map( A1 => n162, A2 => n815, B => n453, C 
                           => n454, Y => crossbar_out(367));
   U659 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(175), A2 => n155, 
                           B1 => crossbar_in(303), B2 => n150, C1 => 
                           crossbar_in(239), C2 => n145, Y => n454);
   U660 : OAI211xp5_ASAP7_75t_R port map( A1 => n162, A2 => n816, B => n455, C 
                           => n456, Y => crossbar_out(366));
   U661 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(174), A2 => n155, 
                           B1 => crossbar_in(302), B2 => n150, C1 => 
                           crossbar_in(238), C2 => n145, Y => n456);
   U662 : OAI211xp5_ASAP7_75t_R port map( A1 => n162, A2 => n817, B => n457, C 
                           => n458, Y => crossbar_out(365));
   U663 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(173), A2 => n155, 
                           B1 => crossbar_in(301), B2 => n150, C1 => 
                           crossbar_in(237), C2 => n145, Y => n458);
   U664 : OAI211xp5_ASAP7_75t_R port map( A1 => n161, A2 => n818, B => n459, C 
                           => n460, Y => crossbar_out(364));
   U665 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(172), A2 => n155, 
                           B1 => crossbar_in(300), B2 => n150, C1 => 
                           crossbar_in(236), C2 => n145, Y => n460);
   U666 : OAI211xp5_ASAP7_75t_R port map( A1 => n161, A2 => n819, B => n461, C 
                           => n462, Y => crossbar_out(363));
   U667 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(171), A2 => n156, 
                           B1 => crossbar_in(299), B2 => n151, C1 => 
                           crossbar_in(235), C2 => n146, Y => n462);
   U668 : OAI211xp5_ASAP7_75t_R port map( A1 => n161, A2 => n820, B => n463, C 
                           => n464, Y => crossbar_out(362));
   U669 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(170), A2 => n156, 
                           B1 => crossbar_in(298), B2 => n151, C1 => 
                           crossbar_in(234), C2 => n146, Y => n464);
   U670 : OAI211xp5_ASAP7_75t_R port map( A1 => n161, A2 => n821, B => n465, C 
                           => n466, Y => crossbar_out(361));
   U671 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(169), A2 => n156, 
                           B1 => crossbar_in(297), B2 => n151, C1 => 
                           crossbar_in(233), C2 => n146, Y => n466);
   U672 : OAI211xp5_ASAP7_75t_R port map( A1 => n161, A2 => n822, B => n467, C 
                           => n468, Y => crossbar_out(360));
   U673 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(168), A2 => n156, 
                           B1 => crossbar_in(296), B2 => n151, C1 => 
                           crossbar_in(232), C2 => n146, Y => n468);
   U674 : OAI211xp5_ASAP7_75t_R port map( A1 => n161, A2 => n390, B => n469, C 
                           => n470, Y => crossbar_out(323));
   U675 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(131), A2 => n156, 
                           B1 => crossbar_in(259), B2 => n151, C1 => 
                           crossbar_in(195), C2 => n146, Y => n470);
   U676 : OAI211xp5_ASAP7_75t_R port map( A1 => n161, A2 => n823, B => n471, C 
                           => n472, Y => crossbar_out(359));
   U677 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(167), A2 => n156, 
                           B1 => crossbar_in(295), B2 => n151, C1 => 
                           crossbar_in(231), C2 => n146, Y => n472);
   U678 : OAI211xp5_ASAP7_75t_R port map( A1 => n161, A2 => n824, B => n473, C 
                           => n474, Y => crossbar_out(358));
   U679 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(166), A2 => n156, 
                           B1 => crossbar_in(294), B2 => n151, C1 => 
                           crossbar_in(230), C2 => n146, Y => n474);
   U680 : OAI211xp5_ASAP7_75t_R port map( A1 => n161, A2 => n825, B => n475, C 
                           => n476, Y => crossbar_out(357));
   U681 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(165), A2 => n156, 
                           B1 => crossbar_in(293), B2 => n151, C1 => 
                           crossbar_in(229), C2 => n146, Y => n476);
   U682 : OAI211xp5_ASAP7_75t_R port map( A1 => n161, A2 => n826, B => n477, C 
                           => n478, Y => crossbar_out(356));
   U683 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(164), A2 => n156, 
                           B1 => crossbar_in(292), B2 => n151, C1 => 
                           crossbar_in(228), C2 => n146, Y => n478);
   U684 : OAI211xp5_ASAP7_75t_R port map( A1 => n161, A2 => n827, B => n479, C 
                           => n480, Y => crossbar_out(355));
   U685 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(163), A2 => n156, 
                           B1 => crossbar_in(291), B2 => n151, C1 => 
                           crossbar_in(227), C2 => n146, Y => n480);
   U686 : OAI211xp5_ASAP7_75t_R port map( A1 => n161, A2 => n828, B => n481, C 
                           => n482, Y => crossbar_out(354));
   U687 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(162), A2 => n156, 
                           B1 => crossbar_in(290), B2 => n151, C1 => 
                           crossbar_in(226), C2 => n146, Y => n482);
   U688 : OAI211xp5_ASAP7_75t_R port map( A1 => n161, A2 => n829, B => n483, C 
                           => n484, Y => crossbar_out(353));
   U689 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(161), A2 => n156, 
                           B1 => crossbar_in(289), B2 => n151, C1 => 
                           crossbar_in(225), C2 => n146, Y => n484);
   U690 : OAI211xp5_ASAP7_75t_R port map( A1 => n160, A2 => n830, B => n485, C 
                           => n486, Y => crossbar_out(352));
   U691 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(160), A2 => n156, 
                           B1 => crossbar_in(288), B2 => n151, C1 => 
                           crossbar_in(224), C2 => n146, Y => n486);
   U692 : OAI211xp5_ASAP7_75t_R port map( A1 => n160, A2 => n831, B => n487, C 
                           => n488, Y => crossbar_out(351));
   U693 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(159), A2 => n157, 
                           B1 => crossbar_in(287), B2 => n152, C1 => 
                           crossbar_in(223), C2 => n147, Y => n488);
   U694 : OAI211xp5_ASAP7_75t_R port map( A1 => n160, A2 => n832, B => n489, C 
                           => n490, Y => crossbar_out(350));
   U695 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(158), A2 => n157, 
                           B1 => crossbar_in(286), B2 => n152, C1 => 
                           crossbar_in(222), C2 => n147, Y => n490);
   U696 : OAI211xp5_ASAP7_75t_R port map( A1 => n160, A2 => n391, B => n491, C 
                           => n492, Y => crossbar_out(322));
   U697 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(130), A2 => n157, 
                           B1 => crossbar_in(258), B2 => n152, C1 => 
                           crossbar_in(194), C2 => n147, Y => n492);
   U698 : OAI211xp5_ASAP7_75t_R port map( A1 => n160, A2 => n364, B => n493, C 
                           => n494, Y => crossbar_out(349));
   U699 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(157), A2 => n157, 
                           B1 => crossbar_in(285), B2 => n152, C1 => 
                           crossbar_in(221), C2 => n147, Y => n494);
   U700 : OAI211xp5_ASAP7_75t_R port map( A1 => n160, A2 => n365, B => n495, C 
                           => n496, Y => crossbar_out(348));
   U701 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(156), A2 => n157, 
                           B1 => crossbar_in(284), B2 => n152, C1 => 
                           crossbar_in(220), C2 => n147, Y => n496);
   U702 : OAI211xp5_ASAP7_75t_R port map( A1 => n160, A2 => n366, B => n497, C 
                           => n498, Y => crossbar_out(347));
   U703 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(155), A2 => n157, 
                           B1 => crossbar_in(283), B2 => n152, C1 => 
                           crossbar_in(219), C2 => n147, Y => n498);
   U704 : OAI211xp5_ASAP7_75t_R port map( A1 => n160, A2 => n367, B => n499, C 
                           => n500, Y => crossbar_out(346));
   U705 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(154), A2 => n157, 
                           B1 => crossbar_in(282), B2 => n152, C1 => 
                           crossbar_in(218), C2 => n147, Y => n500);
   U706 : OAI211xp5_ASAP7_75t_R port map( A1 => n160, A2 => n368, B => n501, C 
                           => n502, Y => crossbar_out(345));
   U707 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(153), A2 => n157, 
                           B1 => crossbar_in(281), B2 => n152, C1 => 
                           crossbar_in(217), C2 => n147, Y => n502);
   U708 : OAI211xp5_ASAP7_75t_R port map( A1 => n160, A2 => n369, B => n503, C 
                           => n504, Y => crossbar_out(344));
   U709 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(152), A2 => n157, 
                           B1 => crossbar_in(280), B2 => n152, C1 => 
                           crossbar_in(216), C2 => n147, Y => n504);
   U710 : OAI211xp5_ASAP7_75t_R port map( A1 => n160, A2 => n370, B => n505, C 
                           => n506, Y => crossbar_out(343));
   U711 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(151), A2 => n157, 
                           B1 => crossbar_in(279), B2 => n152, C1 => 
                           crossbar_in(215), C2 => n147, Y => n506);
   U712 : OAI211xp5_ASAP7_75t_R port map( A1 => n160, A2 => n371, B => n507, C 
                           => n508, Y => crossbar_out(342));
   U713 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(150), A2 => n157, 
                           B1 => crossbar_in(278), B2 => n152, C1 => 
                           crossbar_in(214), C2 => n147, Y => n508);
   U714 : OAI211xp5_ASAP7_75t_R port map( A1 => n160, A2 => n372, B => n509, C 
                           => n510, Y => crossbar_out(341));
   U715 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(149), A2 => n157, 
                           B1 => crossbar_in(277), B2 => n152, C1 => 
                           crossbar_in(213), C2 => n147, Y => n510);
   U716 : OAI211xp5_ASAP7_75t_R port map( A1 => n159, A2 => n373, B => n511, C 
                           => n512, Y => crossbar_out(340));
   U717 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(148), A2 => n157, 
                           B1 => crossbar_in(276), B2 => n152, C1 => 
                           crossbar_in(212), C2 => n147, Y => n512);
   U718 : OAI211xp5_ASAP7_75t_R port map( A1 => n159, A2 => n392, B => n513, C 
                           => n514, Y => crossbar_out(321));
   U719 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(129), A2 => n158, 
                           B1 => crossbar_in(257), B2 => n153, C1 => 
                           crossbar_in(193), C2 => n148, Y => n514);
   U720 : OAI211xp5_ASAP7_75t_R port map( A1 => n159, A2 => n374, B => n515, C 
                           => n516, Y => crossbar_out(339));
   U721 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(147), A2 => n158, 
                           B1 => crossbar_in(275), B2 => n153, C1 => 
                           crossbar_in(211), C2 => n148, Y => n516);
   U722 : OAI211xp5_ASAP7_75t_R port map( A1 => n159, A2 => n375, B => n517, C 
                           => n518, Y => crossbar_out(338));
   U723 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(146), A2 => n158, 
                           B1 => crossbar_in(274), B2 => n153, C1 => 
                           crossbar_in(210), C2 => n148, Y => n518);
   U724 : OAI211xp5_ASAP7_75t_R port map( A1 => n159, A2 => n376, B => n519, C 
                           => n520, Y => crossbar_out(337));
   U725 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(145), A2 => n158, 
                           B1 => crossbar_in(273), B2 => n153, C1 => 
                           crossbar_in(209), C2 => n148, Y => n520);
   U726 : OAI211xp5_ASAP7_75t_R port map( A1 => n159, A2 => n377, B => n521, C 
                           => n522, Y => crossbar_out(336));
   U727 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(144), A2 => n158, 
                           B1 => crossbar_in(272), B2 => n153, C1 => 
                           crossbar_in(208), C2 => n148, Y => n522);
   U728 : OAI211xp5_ASAP7_75t_R port map( A1 => n159, A2 => n378, B => n523, C 
                           => n524, Y => crossbar_out(335));
   U729 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(143), A2 => n158, 
                           B1 => crossbar_in(271), B2 => n153, C1 => 
                           crossbar_in(207), C2 => n148, Y => n524);
   U730 : OAI211xp5_ASAP7_75t_R port map( A1 => n159, A2 => n379, B => n525, C 
                           => n526, Y => crossbar_out(334));
   U731 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(142), A2 => n158, 
                           B1 => crossbar_in(270), B2 => n153, C1 => 
                           crossbar_in(206), C2 => n148, Y => n526);
   U732 : OAI211xp5_ASAP7_75t_R port map( A1 => n159, A2 => n380, B => n527, C 
                           => n528, Y => crossbar_out(333));
   U733 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(141), A2 => n158, 
                           B1 => crossbar_in(269), B2 => n153, C1 => 
                           crossbar_in(205), C2 => n148, Y => n528);
   U734 : OAI211xp5_ASAP7_75t_R port map( A1 => n159, A2 => n381, B => n529, C 
                           => n530, Y => crossbar_out(332));
   U735 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(140), A2 => n158, 
                           B1 => crossbar_in(268), B2 => n153, C1 => 
                           crossbar_in(204), C2 => n148, Y => n530);
   U736 : OAI211xp5_ASAP7_75t_R port map( A1 => n159, A2 => n382, B => n531, C 
                           => n532, Y => crossbar_out(331));
   U737 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(139), A2 => n158, 
                           B1 => crossbar_in(267), B2 => n153, C1 => 
                           crossbar_in(203), C2 => n148, Y => n532);
   U738 : OAI211xp5_ASAP7_75t_R port map( A1 => n159, A2 => n383, B => n533, C 
                           => n534, Y => crossbar_out(330));
   U739 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(138), A2 => n158, 
                           B1 => crossbar_in(266), B2 => n153, C1 => 
                           crossbar_in(202), C2 => n148, Y => n534);
   U740 : OAI211xp5_ASAP7_75t_R port map( A1 => n159, A2 => n393, B => n535, C 
                           => n536, Y => crossbar_out(320));
   U741 : AOI222xp33_ASAP7_75t_R port map( A1 => crossbar_in(128), A2 => n158, 
                           B1 => crossbar_in(256), B2 => n153, C1 => 
                           crossbar_in(192), C2 => n148, Y => n536);
   U742 : NAND3xp33_ASAP7_75t_R port map( A => n898, B => n897, C => n899, Y =>
                           n403);
   U743 : OAI222xp33_ASAP7_75t_R port map( A1 => n976, A2 => n18, B1 => n320, 
                           B2 => n131, C1 => n853, C2 => n12, Y => 
                           crossbar_out(265));
   U744 : OAI222xp33_ASAP7_75t_R port map( A1 => n975, A2 => n18, B1 => n321, 
                           B2 => n131, C1 => n854, C2 => n12, Y => 
                           crossbar_out(264));
   U745 : OAI222xp33_ASAP7_75t_R port map( A1 => n974, A2 => n18, B1 => n322, 
                           B2 => n131, C1 => n855, C2 => n12, Y => 
                           crossbar_out(263));
   U746 : OAI222xp33_ASAP7_75t_R port map( A1 => n973, A2 => n18, B1 => n323, 
                           B2 => n131, C1 => n856, C2 => n12, Y => 
                           crossbar_out(262));
   U747 : OAI222xp33_ASAP7_75t_R port map( A1 => n972, A2 => n17, B1 => n330, 
                           B2 => n130, C1 => n863, C2 => n11, Y => 
                           crossbar_out(319));
   U748 : OAI222xp33_ASAP7_75t_R port map( A1 => n971, A2 => n17, B1 => n331, 
                           B2 => n130, C1 => n864, C2 => n11, Y => 
                           crossbar_out(318));
   U749 : OAI222xp33_ASAP7_75t_R port map( A1 => n970, A2 => n17, B1 => n332, 
                           B2 => n130, C1 => n865, C2 => n11, Y => 
                           crossbar_out(317));
   U750 : OAI222xp33_ASAP7_75t_R port map( A1 => n969, A2 => n17, B1 => n333, 
                           B2 => n130, C1 => n866, C2 => n11, Y => 
                           crossbar_out(316));
   U751 : OAI222xp33_ASAP7_75t_R port map( A1 => n968, A2 => n17, B1 => n324, 
                           B2 => n130, C1 => n857, C2 => n11, Y => 
                           crossbar_out(261));
   U752 : OAI222xp33_ASAP7_75t_R port map( A1 => n967, A2 => n17, B1 => n334, 
                           B2 => n130, C1 => n867, C2 => n11, Y => 
                           crossbar_out(315));
   U753 : OAI222xp33_ASAP7_75t_R port map( A1 => n966, A2 => n17, B1 => n335, 
                           B2 => n130, C1 => n868, C2 => n11, Y => 
                           crossbar_out(314));
   U754 : OAI222xp33_ASAP7_75t_R port map( A1 => n965, A2 => n17, B1 => n336, 
                           B2 => n130, C1 => n869, C2 => n11, Y => 
                           crossbar_out(313));
   U755 : OAI222xp33_ASAP7_75t_R port map( A1 => n964, A2 => n17, B1 => n337, 
                           B2 => n130, C1 => n870, C2 => n11, Y => 
                           crossbar_out(312));
   U756 : OAI222xp33_ASAP7_75t_R port map( A1 => n963, A2 => n17, B1 => n338, 
                           B2 => n130, C1 => n871, C2 => n11, Y => 
                           crossbar_out(311));
   U757 : OAI222xp33_ASAP7_75t_R port map( A1 => n962, A2 => n17, B1 => n339, 
                           B2 => n130, C1 => n872, C2 => n11, Y => 
                           crossbar_out(310));
   U758 : OAI222xp33_ASAP7_75t_R port map( A1 => n961, A2 => n17, B1 => n340, 
                           B2 => n130, C1 => n873, C2 => n11, Y => 
                           crossbar_out(309));
   U759 : OAI222xp33_ASAP7_75t_R port map( A1 => n960, A2 => n16, B1 => n341, 
                           B2 => n129, C1 => n874, C2 => n10, Y => 
                           crossbar_out(308));
   U760 : OAI222xp33_ASAP7_75t_R port map( A1 => n959, A2 => n16, B1 => n342, 
                           B2 => n129, C1 => n875, C2 => n10, Y => 
                           crossbar_out(307));
   U761 : OAI222xp33_ASAP7_75t_R port map( A1 => n958, A2 => n16, B1 => n343, 
                           B2 => n129, C1 => n876, C2 => n10, Y => 
                           crossbar_out(306));
   U762 : OAI222xp33_ASAP7_75t_R port map( A1 => n957, A2 => n16, B1 => n325, 
                           B2 => n129, C1 => n858, C2 => n10, Y => 
                           crossbar_out(260));
   U763 : OAI222xp33_ASAP7_75t_R port map( A1 => n956, A2 => n16, B1 => n344, 
                           B2 => n129, C1 => n877, C2 => n10, Y => 
                           crossbar_out(305));
   U764 : OAI222xp33_ASAP7_75t_R port map( A1 => n955, A2 => n16, B1 => n345, 
                           B2 => n129, C1 => n878, C2 => n10, Y => 
                           crossbar_out(304));
   U765 : OAI222xp33_ASAP7_75t_R port map( A1 => n954, A2 => n16, B1 => n346, 
                           B2 => n129, C1 => n879, C2 => n10, Y => 
                           crossbar_out(303));
   U766 : OAI222xp33_ASAP7_75t_R port map( A1 => n953, A2 => n16, B1 => n347, 
                           B2 => n129, C1 => n880, C2 => n10, Y => 
                           crossbar_out(302));
   U767 : OAI222xp33_ASAP7_75t_R port map( A1 => n952, A2 => n16, B1 => n348, 
                           B2 => n129, C1 => n881, C2 => n10, Y => 
                           crossbar_out(301));
   U768 : OAI222xp33_ASAP7_75t_R port map( A1 => n951, A2 => n16, B1 => n349, 
                           B2 => n129, C1 => n882, C2 => n10, Y => 
                           crossbar_out(300));
   U769 : OAI222xp33_ASAP7_75t_R port map( A1 => n950, A2 => n16, B1 => n350, 
                           B2 => n129, C1 => n883, C2 => n10, Y => 
                           crossbar_out(299));
   U770 : OAI222xp33_ASAP7_75t_R port map( A1 => n949, A2 => n16, B1 => n351, 
                           B2 => n129, C1 => n884, C2 => n10, Y => 
                           crossbar_out(298));
   U771 : OAI222xp33_ASAP7_75t_R port map( A1 => n948, A2 => n15, B1 => n352, 
                           B2 => n128, C1 => n885, C2 => n9, Y => 
                           crossbar_out(297));
   U772 : OAI222xp33_ASAP7_75t_R port map( A1 => n947, A2 => n15, B1 => n353, 
                           B2 => n128, C1 => n886, C2 => n9, Y => 
                           crossbar_out(296));
   U773 : OAI222xp33_ASAP7_75t_R port map( A1 => n946, A2 => n15, B1 => n326, 
                           B2 => n128, C1 => n859, C2 => n9, Y => 
                           crossbar_out(259));
   U774 : OAI222xp33_ASAP7_75t_R port map( A1 => n945, A2 => n15, B1 => n354, 
                           B2 => n128, C1 => n887, C2 => n9, Y => 
                           crossbar_out(295));
   U775 : OAI222xp33_ASAP7_75t_R port map( A1 => n944, A2 => n15, B1 => n355, 
                           B2 => n128, C1 => n888, C2 => n9, Y => 
                           crossbar_out(294));
   U776 : OAI222xp33_ASAP7_75t_R port map( A1 => n943, A2 => n15, B1 => n356, 
                           B2 => n128, C1 => n889, C2 => n9, Y => 
                           crossbar_out(293));
   U777 : OAI222xp33_ASAP7_75t_R port map( A1 => n942, A2 => n15, B1 => n357, 
                           B2 => n128, C1 => n890, C2 => n9, Y => 
                           crossbar_out(292));
   U778 : OAI222xp33_ASAP7_75t_R port map( A1 => n941, A2 => n15, B1 => n358, 
                           B2 => n128, C1 => n891, C2 => n9, Y => 
                           crossbar_out(291));
   U779 : OAI222xp33_ASAP7_75t_R port map( A1 => n940, A2 => n15, B1 => n359, 
                           B2 => n128, C1 => n892, C2 => n9, Y => 
                           crossbar_out(290));
   U780 : OAI222xp33_ASAP7_75t_R port map( A1 => n939, A2 => n15, B1 => n360, 
                           B2 => n128, C1 => n893, C2 => n9, Y => 
                           crossbar_out(289));
   U781 : OAI222xp33_ASAP7_75t_R port map( A1 => n938, A2 => n15, B1 => n361, 
                           B2 => n128, C1 => n894, C2 => n9, Y => 
                           crossbar_out(288));
   U782 : OAI222xp33_ASAP7_75t_R port map( A1 => n937, A2 => n15, B1 => n362, 
                           B2 => n128, C1 => n895, C2 => n9, Y => 
                           crossbar_out(287));
   U783 : OAI222xp33_ASAP7_75t_R port map( A1 => n936, A2 => n14, B1 => n363, 
                           B2 => n127, C1 => n896, C2 => n8, Y => 
                           crossbar_out(286));
   U784 : OAI222xp33_ASAP7_75t_R port map( A1 => n935, A2 => n14, B1 => n327, 
                           B2 => n127, C1 => n860, C2 => n8, Y => 
                           crossbar_out(258));
   U785 : OAI222xp33_ASAP7_75t_R port map( A1 => n934, A2 => n14, B1 => n300, 
                           B2 => n127, C1 => n833, C2 => n8, Y => 
                           crossbar_out(285));
   U786 : OAI222xp33_ASAP7_75t_R port map( A1 => n933, A2 => n14, B1 => n301, 
                           B2 => n127, C1 => n834, C2 => n8, Y => 
                           crossbar_out(284));
   U787 : OAI222xp33_ASAP7_75t_R port map( A1 => n932, A2 => n14, B1 => n302, 
                           B2 => n127, C1 => n835, C2 => n8, Y => 
                           crossbar_out(283));
   U788 : OAI222xp33_ASAP7_75t_R port map( A1 => n931, A2 => n14, B1 => n303, 
                           B2 => n127, C1 => n836, C2 => n8, Y => 
                           crossbar_out(282));
   U789 : OAI222xp33_ASAP7_75t_R port map( A1 => n930, A2 => n14, B1 => n304, 
                           B2 => n127, C1 => n837, C2 => n8, Y => 
                           crossbar_out(281));
   U790 : OAI222xp33_ASAP7_75t_R port map( A1 => n929, A2 => n14, B1 => n305, 
                           B2 => n127, C1 => n838, C2 => n8, Y => 
                           crossbar_out(280));
   U791 : OAI222xp33_ASAP7_75t_R port map( A1 => n928, A2 => n14, B1 => n306, 
                           B2 => n127, C1 => n839, C2 => n8, Y => 
                           crossbar_out(279));
   U792 : OAI222xp33_ASAP7_75t_R port map( A1 => n927, A2 => n14, B1 => n307, 
                           B2 => n127, C1 => n840, C2 => n8, Y => 
                           crossbar_out(278));
   U793 : OAI222xp33_ASAP7_75t_R port map( A1 => n926, A2 => n14, B1 => n308, 
                           B2 => n127, C1 => n841, C2 => n8, Y => 
                           crossbar_out(277));
   U794 : OAI222xp33_ASAP7_75t_R port map( A1 => n925, A2 => n14, B1 => n309, 
                           B2 => n127, C1 => n842, C2 => n8, Y => 
                           crossbar_out(276));
   U795 : OAI222xp33_ASAP7_75t_R port map( A1 => n924, A2 => n13, B1 => n328, 
                           B2 => n126, C1 => n861, C2 => n7, Y => 
                           crossbar_out(257));
   U796 : OAI222xp33_ASAP7_75t_R port map( A1 => n923, A2 => n13, B1 => n310, 
                           B2 => n126, C1 => n843, C2 => n7, Y => 
                           crossbar_out(275));
   U797 : OAI222xp33_ASAP7_75t_R port map( A1 => n922, A2 => n13, B1 => n311, 
                           B2 => n126, C1 => n844, C2 => n7, Y => 
                           crossbar_out(274));
   U798 : OAI222xp33_ASAP7_75t_R port map( A1 => n921, A2 => n13, B1 => n312, 
                           B2 => n126, C1 => n845, C2 => n7, Y => 
                           crossbar_out(273));
   U799 : OAI222xp33_ASAP7_75t_R port map( A1 => n920, A2 => n13, B1 => n313, 
                           B2 => n126, C1 => n846, C2 => n7, Y => 
                           crossbar_out(272));
   U800 : OAI222xp33_ASAP7_75t_R port map( A1 => n919, A2 => n13, B1 => n314, 
                           B2 => n126, C1 => n847, C2 => n7, Y => 
                           crossbar_out(271));
   U801 : OAI222xp33_ASAP7_75t_R port map( A1 => n918, A2 => n13, B1 => n315, 
                           B2 => n126, C1 => n848, C2 => n7, Y => 
                           crossbar_out(270));
   U802 : OAI222xp33_ASAP7_75t_R port map( A1 => n917, A2 => n13, B1 => n316, 
                           B2 => n126, C1 => n849, C2 => n7, Y => 
                           crossbar_out(269));
   U803 : OAI222xp33_ASAP7_75t_R port map( A1 => n916, A2 => n13, B1 => n317, 
                           B2 => n126, C1 => n850, C2 => n7, Y => 
                           crossbar_out(268));
   U804 : OAI222xp33_ASAP7_75t_R port map( A1 => n915, A2 => n13, B1 => n318, 
                           B2 => n126, C1 => n851, C2 => n7, Y => 
                           crossbar_out(267));
   U805 : OAI222xp33_ASAP7_75t_R port map( A1 => n914, A2 => n13, B1 => n319, 
                           B2 => n126, C1 => n852, C2 => n7, Y => 
                           crossbar_out(266));
   U806 : OAI222xp33_ASAP7_75t_R port map( A1 => n913, A2 => n13, B1 => n329, 
                           B2 => n126, C1 => n862, C2 => n7, Y => 
                           crossbar_out(256));
   U807 : OAI221xp5_ASAP7_75t_R port map( A1 => n256, A2 => n120, B1 => n976, 
                           B2 => n6, C => n539, Y => crossbar_out(201));
   U808 : AOI222xp33_ASAP7_75t_R port map( A1 => n114, A2 => crossbar_in(329), 
                           B1 => n108, B2 => crossbar_in(137), C1 => n102, C2 
                           => crossbar_in(73), Y => n539);
   U809 : OAI221xp5_ASAP7_75t_R port map( A1 => n257, A2 => n120, B1 => n975, 
                           B2 => n6, C => n543, Y => crossbar_out(200));
   U810 : AOI222xp33_ASAP7_75t_R port map( A1 => n114, A2 => crossbar_in(328), 
                           B1 => n108, B2 => crossbar_in(136), C1 => n102, C2 
                           => crossbar_in(72), Y => n543);
   U811 : OAI221xp5_ASAP7_75t_R port map( A1 => n258, A2 => n120, B1 => n974, 
                           B2 => n6, C => n544, Y => crossbar_out(199));
   U812 : AOI222xp33_ASAP7_75t_R port map( A1 => n114, A2 => crossbar_in(327), 
                           B1 => n108, B2 => crossbar_in(135), C1 => n102, C2 
                           => crossbar_in(71), Y => n544);
   U813 : OAI221xp5_ASAP7_75t_R port map( A1 => n259, A2 => n120, B1 => n973, 
                           B2 => n6, C => n545, Y => crossbar_out(198));
   U814 : AOI222xp33_ASAP7_75t_R port map( A1 => n114, A2 => crossbar_in(326), 
                           B1 => n108, B2 => crossbar_in(134), C1 => n102, C2 
                           => crossbar_in(70), Y => n545);
   U815 : OAI221xp5_ASAP7_75t_R port map( A1 => n266, A2 => n120, B1 => n972, 
                           B2 => n5, C => n546, Y => crossbar_out(255));
   U816 : AOI222xp33_ASAP7_75t_R port map( A1 => n114, A2 => crossbar_in(383), 
                           B1 => n108, B2 => crossbar_in(191), C1 => n102, C2 
                           => crossbar_in(127), Y => n546);
   U817 : OAI221xp5_ASAP7_75t_R port map( A1 => n267, A2 => n120, B1 => n971, 
                           B2 => n5, C => n547, Y => crossbar_out(254));
   U818 : AOI222xp33_ASAP7_75t_R port map( A1 => n114, A2 => crossbar_in(382), 
                           B1 => n108, B2 => crossbar_in(190), C1 => n102, C2 
                           => crossbar_in(126), Y => n547);
   U819 : OAI221xp5_ASAP7_75t_R port map( A1 => n268, A2 => n120, B1 => n970, 
                           B2 => n5, C => n548, Y => crossbar_out(253));
   U820 : AOI222xp33_ASAP7_75t_R port map( A1 => n114, A2 => crossbar_in(381), 
                           B1 => n108, B2 => crossbar_in(189), C1 => n102, C2 
                           => crossbar_in(125), Y => n548);
   U821 : OAI221xp5_ASAP7_75t_R port map( A1 => n269, A2 => n120, B1 => n969, 
                           B2 => n5, C => n549, Y => crossbar_out(252));
   U822 : AOI222xp33_ASAP7_75t_R port map( A1 => n114, A2 => crossbar_in(380), 
                           B1 => n108, B2 => crossbar_in(188), C1 => n102, C2 
                           => crossbar_in(124), Y => n549);
   U823 : OAI221xp5_ASAP7_75t_R port map( A1 => n260, A2 => n120, B1 => n968, 
                           B2 => n5, C => n550, Y => crossbar_out(197));
   U824 : AOI222xp33_ASAP7_75t_R port map( A1 => n114, A2 => crossbar_in(325), 
                           B1 => n108, B2 => crossbar_in(133), C1 => n102, C2 
                           => crossbar_in(69), Y => n550);
   U825 : OAI221xp5_ASAP7_75t_R port map( A1 => n270, A2 => n120, B1 => n967, 
                           B2 => n5, C => n551, Y => crossbar_out(251));
   U826 : AOI222xp33_ASAP7_75t_R port map( A1 => n114, A2 => crossbar_in(379), 
                           B1 => n108, B2 => crossbar_in(187), C1 => n102, C2 
                           => crossbar_in(123), Y => n551);
   U827 : OAI221xp5_ASAP7_75t_R port map( A1 => n271, A2 => n120, B1 => n966, 
                           B2 => n5, C => n552, Y => crossbar_out(250));
   U828 : AOI222xp33_ASAP7_75t_R port map( A1 => n114, A2 => crossbar_in(378), 
                           B1 => n108, B2 => crossbar_in(186), C1 => n102, C2 
                           => crossbar_in(122), Y => n552);
   U829 : OAI221xp5_ASAP7_75t_R port map( A1 => n272, A2 => n120, B1 => n965, 
                           B2 => n5, C => n553, Y => crossbar_out(249));
   U830 : AOI222xp33_ASAP7_75t_R port map( A1 => n114, A2 => crossbar_in(377), 
                           B1 => n108, B2 => crossbar_in(185), C1 => n102, C2 
                           => crossbar_in(121), Y => n553);
   U831 : OAI221xp5_ASAP7_75t_R port map( A1 => n273, A2 => n121, B1 => n964, 
                           B2 => n5, C => n554, Y => crossbar_out(248));
   U832 : AOI222xp33_ASAP7_75t_R port map( A1 => n115, A2 => crossbar_in(376), 
                           B1 => n109, B2 => crossbar_in(184), C1 => n103, C2 
                           => crossbar_in(120), Y => n554);
   U833 : OAI221xp5_ASAP7_75t_R port map( A1 => n274, A2 => n121, B1 => n963, 
                           B2 => n5, C => n555, Y => crossbar_out(247));
   U834 : AOI222xp33_ASAP7_75t_R port map( A1 => n115, A2 => crossbar_in(375), 
                           B1 => n109, B2 => crossbar_in(183), C1 => n103, C2 
                           => crossbar_in(119), Y => n555);
   U835 : OAI221xp5_ASAP7_75t_R port map( A1 => n275, A2 => n121, B1 => n962, 
                           B2 => n5, C => n556, Y => crossbar_out(246));
   U836 : AOI222xp33_ASAP7_75t_R port map( A1 => n115, A2 => crossbar_in(374), 
                           B1 => n109, B2 => crossbar_in(182), C1 => n103, C2 
                           => crossbar_in(118), Y => n556);
   U837 : OAI221xp5_ASAP7_75t_R port map( A1 => n276, A2 => n121, B1 => n961, 
                           B2 => n5, C => n557, Y => crossbar_out(245));
   U838 : AOI222xp33_ASAP7_75t_R port map( A1 => n115, A2 => crossbar_in(373), 
                           B1 => n109, B2 => crossbar_in(181), C1 => n103, C2 
                           => crossbar_in(117), Y => n557);
   U839 : OAI221xp5_ASAP7_75t_R port map( A1 => n277, A2 => n121, B1 => n960, 
                           B2 => n4, C => n558, Y => crossbar_out(244));
   U840 : AOI222xp33_ASAP7_75t_R port map( A1 => n115, A2 => crossbar_in(372), 
                           B1 => n109, B2 => crossbar_in(180), C1 => n103, C2 
                           => crossbar_in(116), Y => n558);
   U841 : OAI221xp5_ASAP7_75t_R port map( A1 => n278, A2 => n121, B1 => n959, 
                           B2 => n4, C => n559, Y => crossbar_out(243));
   U842 : AOI222xp33_ASAP7_75t_R port map( A1 => n115, A2 => crossbar_in(371), 
                           B1 => n109, B2 => crossbar_in(179), C1 => n103, C2 
                           => crossbar_in(115), Y => n559);
   U843 : OAI221xp5_ASAP7_75t_R port map( A1 => n279, A2 => n121, B1 => n958, 
                           B2 => n4, C => n560, Y => crossbar_out(242));
   U844 : AOI222xp33_ASAP7_75t_R port map( A1 => n115, A2 => crossbar_in(370), 
                           B1 => n109, B2 => crossbar_in(178), C1 => n103, C2 
                           => crossbar_in(114), Y => n560);
   U845 : OAI221xp5_ASAP7_75t_R port map( A1 => n261, A2 => n121, B1 => n957, 
                           B2 => n4, C => n561, Y => crossbar_out(196));
   U846 : AOI222xp33_ASAP7_75t_R port map( A1 => n115, A2 => crossbar_in(324), 
                           B1 => n109, B2 => crossbar_in(132), C1 => n103, C2 
                           => crossbar_in(68), Y => n561);
   U847 : OAI221xp5_ASAP7_75t_R port map( A1 => n280, A2 => n121, B1 => n956, 
                           B2 => n4, C => n562, Y => crossbar_out(241));
   U848 : AOI222xp33_ASAP7_75t_R port map( A1 => n115, A2 => crossbar_in(369), 
                           B1 => n109, B2 => crossbar_in(177), C1 => n103, C2 
                           => crossbar_in(113), Y => n562);
   U849 : OAI221xp5_ASAP7_75t_R port map( A1 => n281, A2 => n121, B1 => n955, 
                           B2 => n4, C => n563, Y => crossbar_out(240));
   U850 : AOI222xp33_ASAP7_75t_R port map( A1 => n115, A2 => crossbar_in(368), 
                           B1 => n109, B2 => crossbar_in(176), C1 => n103, C2 
                           => crossbar_in(112), Y => n563);
   U851 : OAI221xp5_ASAP7_75t_R port map( A1 => n282, A2 => n121, B1 => n954, 
                           B2 => n4, C => n564, Y => crossbar_out(239));
   U852 : AOI222xp33_ASAP7_75t_R port map( A1 => n115, A2 => crossbar_in(367), 
                           B1 => n109, B2 => crossbar_in(175), C1 => n103, C2 
                           => crossbar_in(111), Y => n564);
   U853 : OAI221xp5_ASAP7_75t_R port map( A1 => n283, A2 => n121, B1 => n953, 
                           B2 => n4, C => n565, Y => crossbar_out(238));
   U854 : AOI222xp33_ASAP7_75t_R port map( A1 => n115, A2 => crossbar_in(366), 
                           B1 => n109, B2 => crossbar_in(174), C1 => n103, C2 
                           => crossbar_in(110), Y => n565);
   U855 : OAI221xp5_ASAP7_75t_R port map( A1 => n284, A2 => n122, B1 => n952, 
                           B2 => n4, C => n566, Y => crossbar_out(237));
   U856 : AOI222xp33_ASAP7_75t_R port map( A1 => n116, A2 => crossbar_in(365), 
                           B1 => n110, B2 => crossbar_in(173), C1 => n104, C2 
                           => crossbar_in(109), Y => n566);
   U857 : OAI221xp5_ASAP7_75t_R port map( A1 => n285, A2 => n122, B1 => n951, 
                           B2 => n4, C => n567, Y => crossbar_out(236));
   U858 : AOI222xp33_ASAP7_75t_R port map( A1 => n116, A2 => crossbar_in(364), 
                           B1 => n110, B2 => crossbar_in(172), C1 => n104, C2 
                           => crossbar_in(108), Y => n567);
   U859 : OAI221xp5_ASAP7_75t_R port map( A1 => n286, A2 => n122, B1 => n950, 
                           B2 => n4, C => n568, Y => crossbar_out(235));
   U860 : AOI222xp33_ASAP7_75t_R port map( A1 => n116, A2 => crossbar_in(363), 
                           B1 => n110, B2 => crossbar_in(171), C1 => n104, C2 
                           => crossbar_in(107), Y => n568);
   U861 : OAI221xp5_ASAP7_75t_R port map( A1 => n287, A2 => n122, B1 => n949, 
                           B2 => n4, C => n569, Y => crossbar_out(234));
   U862 : AOI222xp33_ASAP7_75t_R port map( A1 => n116, A2 => crossbar_in(362), 
                           B1 => n110, B2 => crossbar_in(170), C1 => n104, C2 
                           => crossbar_in(106), Y => n569);
   U863 : OAI221xp5_ASAP7_75t_R port map( A1 => n288, A2 => n122, B1 => n948, 
                           B2 => n3, C => n570, Y => crossbar_out(233));
   U864 : AOI222xp33_ASAP7_75t_R port map( A1 => n116, A2 => crossbar_in(361), 
                           B1 => n110, B2 => crossbar_in(169), C1 => n104, C2 
                           => crossbar_in(105), Y => n570);
   U865 : OAI221xp5_ASAP7_75t_R port map( A1 => n289, A2 => n122, B1 => n947, 
                           B2 => n3, C => n571, Y => crossbar_out(232));
   U866 : AOI222xp33_ASAP7_75t_R port map( A1 => n116, A2 => crossbar_in(360), 
                           B1 => n110, B2 => crossbar_in(168), C1 => n104, C2 
                           => crossbar_in(104), Y => n571);
   U867 : OAI221xp5_ASAP7_75t_R port map( A1 => n262, A2 => n122, B1 => n946, 
                           B2 => n3, C => n572, Y => crossbar_out(195));
   U868 : AOI222xp33_ASAP7_75t_R port map( A1 => n116, A2 => crossbar_in(323), 
                           B1 => n110, B2 => crossbar_in(131), C1 => n104, C2 
                           => crossbar_in(67), Y => n572);
   U869 : OAI221xp5_ASAP7_75t_R port map( A1 => n290, A2 => n122, B1 => n945, 
                           B2 => n3, C => n573, Y => crossbar_out(231));
   U870 : AOI222xp33_ASAP7_75t_R port map( A1 => n116, A2 => crossbar_in(359), 
                           B1 => n110, B2 => crossbar_in(167), C1 => n104, C2 
                           => crossbar_in(103), Y => n573);
   U871 : OAI221xp5_ASAP7_75t_R port map( A1 => n291, A2 => n122, B1 => n944, 
                           B2 => n3, C => n574, Y => crossbar_out(230));
   U872 : AOI222xp33_ASAP7_75t_R port map( A1 => n116, A2 => crossbar_in(358), 
                           B1 => n110, B2 => crossbar_in(166), C1 => n104, C2 
                           => crossbar_in(102), Y => n574);
   U873 : OAI221xp5_ASAP7_75t_R port map( A1 => n292, A2 => n122, B1 => n943, 
                           B2 => n3, C => n575, Y => crossbar_out(229));
   U874 : AOI222xp33_ASAP7_75t_R port map( A1 => n116, A2 => crossbar_in(357), 
                           B1 => n110, B2 => crossbar_in(165), C1 => n104, C2 
                           => crossbar_in(101), Y => n575);
   U875 : OAI221xp5_ASAP7_75t_R port map( A1 => n293, A2 => n122, B1 => n942, 
                           B2 => n3, C => n576, Y => crossbar_out(228));
   U876 : AOI222xp33_ASAP7_75t_R port map( A1 => n116, A2 => crossbar_in(356), 
                           B1 => n110, B2 => crossbar_in(164), C1 => n104, C2 
                           => crossbar_in(100), Y => n576);
   U877 : OAI221xp5_ASAP7_75t_R port map( A1 => n294, A2 => n122, B1 => n941, 
                           B2 => n3, C => n577, Y => crossbar_out(227));
   U878 : AOI222xp33_ASAP7_75t_R port map( A1 => n116, A2 => crossbar_in(355), 
                           B1 => n110, B2 => crossbar_in(163), C1 => n104, C2 
                           => crossbar_in(99), Y => n577);
   U879 : OAI221xp5_ASAP7_75t_R port map( A1 => n295, A2 => n123, B1 => n940, 
                           B2 => n3, C => n578, Y => crossbar_out(226));
   U880 : AOI222xp33_ASAP7_75t_R port map( A1 => n117, A2 => crossbar_in(354), 
                           B1 => n111, B2 => crossbar_in(162), C1 => n105, C2 
                           => crossbar_in(98), Y => n578);
   U881 : OAI221xp5_ASAP7_75t_R port map( A1 => n296, A2 => n123, B1 => n939, 
                           B2 => n3, C => n579, Y => crossbar_out(225));
   U882 : AOI222xp33_ASAP7_75t_R port map( A1 => n117, A2 => crossbar_in(353), 
                           B1 => n111, B2 => crossbar_in(161), C1 => n105, C2 
                           => crossbar_in(97), Y => n579);
   U883 : OAI221xp5_ASAP7_75t_R port map( A1 => n297, A2 => n123, B1 => n938, 
                           B2 => n3, C => n580, Y => crossbar_out(224));
   U884 : AOI222xp33_ASAP7_75t_R port map( A1 => n117, A2 => crossbar_in(352), 
                           B1 => n111, B2 => crossbar_in(160), C1 => n105, C2 
                           => crossbar_in(96), Y => n580);
   U885 : OAI221xp5_ASAP7_75t_R port map( A1 => n298, A2 => n123, B1 => n937, 
                           B2 => n3, C => n581, Y => crossbar_out(223));
   U886 : AOI222xp33_ASAP7_75t_R port map( A1 => n117, A2 => crossbar_in(351), 
                           B1 => n111, B2 => crossbar_in(159), C1 => n105, C2 
                           => crossbar_in(95), Y => n581);
   U887 : OAI221xp5_ASAP7_75t_R port map( A1 => n299, A2 => n123, B1 => n936, 
                           B2 => n2, C => n582, Y => crossbar_out(222));
   U888 : AOI222xp33_ASAP7_75t_R port map( A1 => n117, A2 => crossbar_in(350), 
                           B1 => n111, B2 => crossbar_in(158), C1 => n105, C2 
                           => crossbar_in(94), Y => n582);
   U889 : OAI221xp5_ASAP7_75t_R port map( A1 => n263, A2 => n123, B1 => n935, 
                           B2 => n2, C => n583, Y => crossbar_out(194));
   U890 : AOI222xp33_ASAP7_75t_R port map( A1 => n117, A2 => crossbar_in(322), 
                           B1 => n111, B2 => crossbar_in(130), C1 => n105, C2 
                           => crossbar_in(66), Y => n583);
   U891 : OAI221xp5_ASAP7_75t_R port map( A1 => n236, A2 => n123, B1 => n934, 
                           B2 => n2, C => n584, Y => crossbar_out(221));
   U892 : AOI222xp33_ASAP7_75t_R port map( A1 => n117, A2 => crossbar_in(349), 
                           B1 => n111, B2 => crossbar_in(157), C1 => n105, C2 
                           => crossbar_in(93), Y => n584);
   U893 : OAI221xp5_ASAP7_75t_R port map( A1 => n237, A2 => n123, B1 => n933, 
                           B2 => n2, C => n585, Y => crossbar_out(220));
   U894 : AOI222xp33_ASAP7_75t_R port map( A1 => n117, A2 => crossbar_in(348), 
                           B1 => n111, B2 => crossbar_in(156), C1 => n105, C2 
                           => crossbar_in(92), Y => n585);
   U895 : OAI221xp5_ASAP7_75t_R port map( A1 => n238, A2 => n123, B1 => n932, 
                           B2 => n2, C => n586, Y => crossbar_out(219));
   U896 : AOI222xp33_ASAP7_75t_R port map( A1 => n117, A2 => crossbar_in(347), 
                           B1 => n111, B2 => crossbar_in(155), C1 => n105, C2 
                           => crossbar_in(91), Y => n586);
   U897 : OAI221xp5_ASAP7_75t_R port map( A1 => n239, A2 => n123, B1 => n931, 
                           B2 => n2, C => n587, Y => crossbar_out(218));
   U898 : AOI222xp33_ASAP7_75t_R port map( A1 => n117, A2 => crossbar_in(346), 
                           B1 => n111, B2 => crossbar_in(154), C1 => n105, C2 
                           => crossbar_in(90), Y => n587);
   U899 : OAI221xp5_ASAP7_75t_R port map( A1 => n240, A2 => n123, B1 => n930, 
                           B2 => n2, C => n588, Y => crossbar_out(217));
   U900 : AOI222xp33_ASAP7_75t_R port map( A1 => n117, A2 => crossbar_in(345), 
                           B1 => n111, B2 => crossbar_in(153), C1 => n105, C2 
                           => crossbar_in(89), Y => n588);
   U901 : OAI221xp5_ASAP7_75t_R port map( A1 => n241, A2 => n123, B1 => n929, 
                           B2 => n2, C => n589, Y => crossbar_out(216));
   U902 : AOI222xp33_ASAP7_75t_R port map( A1 => n117, A2 => crossbar_in(344), 
                           B1 => n111, B2 => crossbar_in(152), C1 => n105, C2 
                           => crossbar_in(88), Y => n589);
   U903 : OAI221xp5_ASAP7_75t_R port map( A1 => n242, A2 => n124, B1 => n928, 
                           B2 => n2, C => n590, Y => crossbar_out(215));
   U904 : AOI222xp33_ASAP7_75t_R port map( A1 => n118, A2 => crossbar_in(343), 
                           B1 => n112, B2 => crossbar_in(151), C1 => n106, C2 
                           => crossbar_in(87), Y => n590);
   U905 : OAI221xp5_ASAP7_75t_R port map( A1 => n243, A2 => n124, B1 => n927, 
                           B2 => n2, C => n591, Y => crossbar_out(214));
   U906 : AOI222xp33_ASAP7_75t_R port map( A1 => n118, A2 => crossbar_in(342), 
                           B1 => n112, B2 => crossbar_in(150), C1 => n106, C2 
                           => crossbar_in(86), Y => n591);
   U907 : OAI221xp5_ASAP7_75t_R port map( A1 => n244, A2 => n124, B1 => n926, 
                           B2 => n2, C => n592, Y => crossbar_out(213));
   U908 : AOI222xp33_ASAP7_75t_R port map( A1 => n118, A2 => crossbar_in(341), 
                           B1 => n112, B2 => crossbar_in(149), C1 => n106, C2 
                           => crossbar_in(85), Y => n592);
   U909 : OAI221xp5_ASAP7_75t_R port map( A1 => n245, A2 => n124, B1 => n925, 
                           B2 => n2, C => n593, Y => crossbar_out(212));
   U910 : AOI222xp33_ASAP7_75t_R port map( A1 => n118, A2 => crossbar_in(340), 
                           B1 => n112, B2 => crossbar_in(148), C1 => n106, C2 
                           => crossbar_in(84), Y => n593);
   U911 : OAI221xp5_ASAP7_75t_R port map( A1 => n264, A2 => n124, B1 => n924, 
                           B2 => n1, C => n594, Y => crossbar_out(193));
   U912 : AOI222xp33_ASAP7_75t_R port map( A1 => n118, A2 => crossbar_in(321), 
                           B1 => n112, B2 => crossbar_in(129), C1 => n106, C2 
                           => crossbar_in(65), Y => n594);
   U913 : OAI221xp5_ASAP7_75t_R port map( A1 => n246, A2 => n124, B1 => n923, 
                           B2 => n1, C => n595, Y => crossbar_out(211));
   U914 : AOI222xp33_ASAP7_75t_R port map( A1 => n118, A2 => crossbar_in(339), 
                           B1 => n112, B2 => crossbar_in(147), C1 => n106, C2 
                           => crossbar_in(83), Y => n595);
   U915 : OAI221xp5_ASAP7_75t_R port map( A1 => n247, A2 => n124, B1 => n922, 
                           B2 => n1, C => n596, Y => crossbar_out(210));
   U916 : AOI222xp33_ASAP7_75t_R port map( A1 => n118, A2 => crossbar_in(338), 
                           B1 => n112, B2 => crossbar_in(146), C1 => n106, C2 
                           => crossbar_in(82), Y => n596);
   U917 : OAI221xp5_ASAP7_75t_R port map( A1 => n248, A2 => n124, B1 => n921, 
                           B2 => n1, C => n597, Y => crossbar_out(209));
   U918 : AOI222xp33_ASAP7_75t_R port map( A1 => n118, A2 => crossbar_in(337), 
                           B1 => n112, B2 => crossbar_in(145), C1 => n106, C2 
                           => crossbar_in(81), Y => n597);
   U919 : OAI221xp5_ASAP7_75t_R port map( A1 => n249, A2 => n124, B1 => n920, 
                           B2 => n1, C => n598, Y => crossbar_out(208));
   U920 : AOI222xp33_ASAP7_75t_R port map( A1 => n118, A2 => crossbar_in(336), 
                           B1 => n112, B2 => crossbar_in(144), C1 => n106, C2 
                           => crossbar_in(80), Y => n598);
   U921 : OAI221xp5_ASAP7_75t_R port map( A1 => n250, A2 => n124, B1 => n919, 
                           B2 => n1, C => n599, Y => crossbar_out(207));
   U922 : AOI222xp33_ASAP7_75t_R port map( A1 => n118, A2 => crossbar_in(335), 
                           B1 => n112, B2 => crossbar_in(143), C1 => n106, C2 
                           => crossbar_in(79), Y => n599);
   U923 : OAI221xp5_ASAP7_75t_R port map( A1 => n251, A2 => n124, B1 => n918, 
                           B2 => n1, C => n600, Y => crossbar_out(206));
   U924 : AOI222xp33_ASAP7_75t_R port map( A1 => n118, A2 => crossbar_in(334), 
                           B1 => n112, B2 => crossbar_in(142), C1 => n106, C2 
                           => crossbar_in(78), Y => n600);
   U925 : OAI221xp5_ASAP7_75t_R port map( A1 => n252, A2 => n124, B1 => n917, 
                           B2 => n1, C => n601, Y => crossbar_out(205));
   U926 : AOI222xp33_ASAP7_75t_R port map( A1 => n118, A2 => crossbar_in(333), 
                           B1 => n112, B2 => crossbar_in(141), C1 => n106, C2 
                           => crossbar_in(77), Y => n601);
   U927 : OAI221xp5_ASAP7_75t_R port map( A1 => n253, A2 => n125, B1 => n916, 
                           B2 => n1, C => n602, Y => crossbar_out(204));
   U928 : AOI222xp33_ASAP7_75t_R port map( A1 => n119, A2 => crossbar_in(332), 
                           B1 => n113, B2 => crossbar_in(140), C1 => n107, C2 
                           => crossbar_in(76), Y => n602);
   U929 : OAI221xp5_ASAP7_75t_R port map( A1 => n254, A2 => n125, B1 => n915, 
                           B2 => n1, C => n603, Y => crossbar_out(203));
   U930 : AOI222xp33_ASAP7_75t_R port map( A1 => n119, A2 => crossbar_in(331), 
                           B1 => n113, B2 => crossbar_in(139), C1 => n107, C2 
                           => crossbar_in(75), Y => n603);
   U931 : OAI221xp5_ASAP7_75t_R port map( A1 => n255, A2 => n125, B1 => n914, 
                           B2 => n1, C => n604, Y => crossbar_out(202));
   U932 : AOI222xp33_ASAP7_75t_R port map( A1 => n119, A2 => crossbar_in(330), 
                           B1 => n113, B2 => crossbar_in(138), C1 => n107, C2 
                           => crossbar_in(74), Y => n604);
   U933 : OAI221xp5_ASAP7_75t_R port map( A1 => n265, A2 => n125, B1 => n913, 
                           B2 => n1, C => n605, Y => crossbar_out(192));
   U934 : AOI222xp33_ASAP7_75t_R port map( A1 => n119, A2 => crossbar_in(320), 
                           B1 => n113, B2 => crossbar_in(128), C1 => n107, C2 
                           => crossbar_in(64), Y => n605);
   U935 : OAI222xp33_ASAP7_75t_R port map( A1 => n320, A2 => n30, B1 => n256, 
                           B2 => n42, C1 => n976, C2 => n36, Y => 
                           crossbar_out(137));
   U936 : OAI222xp33_ASAP7_75t_R port map( A1 => n321, A2 => n30, B1 => n257, 
                           B2 => n42, C1 => n975, C2 => n36, Y => 
                           crossbar_out(136));
   U937 : OAI222xp33_ASAP7_75t_R port map( A1 => n322, A2 => n30, B1 => n258, 
                           B2 => n42, C1 => n974, C2 => n36, Y => 
                           crossbar_out(135));
   U938 : OAI222xp33_ASAP7_75t_R port map( A1 => n323, A2 => n30, B1 => n259, 
                           B2 => n42, C1 => n973, C2 => n36, Y => 
                           crossbar_out(134));
   U939 : OAI222xp33_ASAP7_75t_R port map( A1 => n330, A2 => n29, B1 => n266, 
                           B2 => n41, C1 => n972, C2 => n35, Y => 
                           crossbar_out(191));
   U940 : OAI222xp33_ASAP7_75t_R port map( A1 => n331, A2 => n29, B1 => n267, 
                           B2 => n41, C1 => n971, C2 => n35, Y => 
                           crossbar_out(190));
   U941 : OAI222xp33_ASAP7_75t_R port map( A1 => n332, A2 => n29, B1 => n268, 
                           B2 => n41, C1 => n970, C2 => n35, Y => 
                           crossbar_out(189));
   U942 : OAI222xp33_ASAP7_75t_R port map( A1 => n333, A2 => n29, B1 => n269, 
                           B2 => n41, C1 => n969, C2 => n35, Y => 
                           crossbar_out(188));
   U943 : OAI222xp33_ASAP7_75t_R port map( A1 => n324, A2 => n29, B1 => n260, 
                           B2 => n41, C1 => n968, C2 => n35, Y => 
                           crossbar_out(133));
   U944 : OAI222xp33_ASAP7_75t_R port map( A1 => n334, A2 => n29, B1 => n270, 
                           B2 => n41, C1 => n967, C2 => n35, Y => 
                           crossbar_out(187));
   U945 : OAI222xp33_ASAP7_75t_R port map( A1 => n335, A2 => n29, B1 => n271, 
                           B2 => n41, C1 => n966, C2 => n35, Y => 
                           crossbar_out(186));
   U946 : OAI222xp33_ASAP7_75t_R port map( A1 => n336, A2 => n29, B1 => n272, 
                           B2 => n41, C1 => n965, C2 => n35, Y => 
                           crossbar_out(185));
   U947 : OAI222xp33_ASAP7_75t_R port map( A1 => n337, A2 => n29, B1 => n273, 
                           B2 => n41, C1 => n964, C2 => n35, Y => 
                           crossbar_out(184));
   U948 : OAI222xp33_ASAP7_75t_R port map( A1 => n338, A2 => n29, B1 => n274, 
                           B2 => n41, C1 => n963, C2 => n35, Y => 
                           crossbar_out(183));
   U949 : OAI222xp33_ASAP7_75t_R port map( A1 => n339, A2 => n29, B1 => n275, 
                           B2 => n41, C1 => n962, C2 => n35, Y => 
                           crossbar_out(182));
   U950 : OAI222xp33_ASAP7_75t_R port map( A1 => n340, A2 => n29, B1 => n276, 
                           B2 => n41, C1 => n961, C2 => n35, Y => 
                           crossbar_out(181));
   U951 : OAI222xp33_ASAP7_75t_R port map( A1 => n341, A2 => n28, B1 => n277, 
                           B2 => n40, C1 => n960, C2 => n34, Y => 
                           crossbar_out(180));
   U952 : OAI222xp33_ASAP7_75t_R port map( A1 => n342, A2 => n28, B1 => n278, 
                           B2 => n40, C1 => n959, C2 => n34, Y => 
                           crossbar_out(179));
   U953 : OAI222xp33_ASAP7_75t_R port map( A1 => n343, A2 => n28, B1 => n279, 
                           B2 => n40, C1 => n958, C2 => n34, Y => 
                           crossbar_out(178));
   U954 : OAI222xp33_ASAP7_75t_R port map( A1 => n325, A2 => n28, B1 => n261, 
                           B2 => n40, C1 => n957, C2 => n34, Y => 
                           crossbar_out(132));
   U955 : OAI222xp33_ASAP7_75t_R port map( A1 => n344, A2 => n28, B1 => n280, 
                           B2 => n40, C1 => n956, C2 => n34, Y => 
                           crossbar_out(177));
   U956 : OAI222xp33_ASAP7_75t_R port map( A1 => n345, A2 => n28, B1 => n281, 
                           B2 => n40, C1 => n955, C2 => n34, Y => 
                           crossbar_out(176));
   U957 : OAI222xp33_ASAP7_75t_R port map( A1 => n346, A2 => n28, B1 => n282, 
                           B2 => n40, C1 => n954, C2 => n34, Y => 
                           crossbar_out(175));
   U958 : OAI222xp33_ASAP7_75t_R port map( A1 => n347, A2 => n28, B1 => n283, 
                           B2 => n40, C1 => n953, C2 => n34, Y => 
                           crossbar_out(174));
   U959 : OAI222xp33_ASAP7_75t_R port map( A1 => n348, A2 => n28, B1 => n284, 
                           B2 => n40, C1 => n952, C2 => n34, Y => 
                           crossbar_out(173));
   U960 : OAI222xp33_ASAP7_75t_R port map( A1 => n349, A2 => n28, B1 => n285, 
                           B2 => n40, C1 => n951, C2 => n34, Y => 
                           crossbar_out(172));
   U961 : OAI222xp33_ASAP7_75t_R port map( A1 => n350, A2 => n28, B1 => n286, 
                           B2 => n40, C1 => n950, C2 => n34, Y => 
                           crossbar_out(171));
   U962 : OAI222xp33_ASAP7_75t_R port map( A1 => n351, A2 => n28, B1 => n287, 
                           B2 => n40, C1 => n949, C2 => n34, Y => 
                           crossbar_out(170));
   U963 : OAI222xp33_ASAP7_75t_R port map( A1 => n352, A2 => n27, B1 => n288, 
                           B2 => n39, C1 => n948, C2 => n33, Y => 
                           crossbar_out(169));
   U964 : OAI222xp33_ASAP7_75t_R port map( A1 => n353, A2 => n27, B1 => n289, 
                           B2 => n39, C1 => n947, C2 => n33, Y => 
                           crossbar_out(168));
   U965 : OAI222xp33_ASAP7_75t_R port map( A1 => n326, A2 => n27, B1 => n262, 
                           B2 => n39, C1 => n946, C2 => n33, Y => 
                           crossbar_out(131));
   U966 : OAI222xp33_ASAP7_75t_R port map( A1 => n354, A2 => n27, B1 => n290, 
                           B2 => n39, C1 => n945, C2 => n33, Y => 
                           crossbar_out(167));
   U967 : OAI222xp33_ASAP7_75t_R port map( A1 => n355, A2 => n27, B1 => n291, 
                           B2 => n39, C1 => n944, C2 => n33, Y => 
                           crossbar_out(166));
   U968 : OAI222xp33_ASAP7_75t_R port map( A1 => n356, A2 => n27, B1 => n292, 
                           B2 => n39, C1 => n943, C2 => n33, Y => 
                           crossbar_out(165));
   U969 : OAI222xp33_ASAP7_75t_R port map( A1 => n357, A2 => n27, B1 => n293, 
                           B2 => n39, C1 => n942, C2 => n33, Y => 
                           crossbar_out(164));
   U970 : OAI222xp33_ASAP7_75t_R port map( A1 => n358, A2 => n27, B1 => n294, 
                           B2 => n39, C1 => n941, C2 => n33, Y => 
                           crossbar_out(163));
   U971 : OAI222xp33_ASAP7_75t_R port map( A1 => n359, A2 => n27, B1 => n295, 
                           B2 => n39, C1 => n940, C2 => n33, Y => 
                           crossbar_out(162));
   U972 : OAI222xp33_ASAP7_75t_R port map( A1 => n360, A2 => n27, B1 => n296, 
                           B2 => n39, C1 => n939, C2 => n33, Y => 
                           crossbar_out(161));
   U973 : OAI222xp33_ASAP7_75t_R port map( A1 => n361, A2 => n27, B1 => n297, 
                           B2 => n39, C1 => n938, C2 => n33, Y => 
                           crossbar_out(160));
   U974 : OAI222xp33_ASAP7_75t_R port map( A1 => n362, A2 => n27, B1 => n298, 
                           B2 => n39, C1 => n937, C2 => n33, Y => 
                           crossbar_out(159));
   U975 : OAI222xp33_ASAP7_75t_R port map( A1 => n363, A2 => n26, B1 => n299, 
                           B2 => n38, C1 => n936, C2 => n32, Y => 
                           crossbar_out(158));
   U976 : OAI222xp33_ASAP7_75t_R port map( A1 => n327, A2 => n26, B1 => n263, 
                           B2 => n38, C1 => n935, C2 => n32, Y => 
                           crossbar_out(130));
   U977 : OAI222xp33_ASAP7_75t_R port map( A1 => n300, A2 => n26, B1 => n236, 
                           B2 => n38, C1 => n934, C2 => n32, Y => 
                           crossbar_out(157));
   U978 : OAI222xp33_ASAP7_75t_R port map( A1 => n301, A2 => n26, B1 => n237, 
                           B2 => n38, C1 => n933, C2 => n32, Y => 
                           crossbar_out(156));
   U979 : OAI222xp33_ASAP7_75t_R port map( A1 => n302, A2 => n26, B1 => n238, 
                           B2 => n38, C1 => n932, C2 => n32, Y => 
                           crossbar_out(155));
   U980 : OAI222xp33_ASAP7_75t_R port map( A1 => n303, A2 => n26, B1 => n239, 
                           B2 => n38, C1 => n931, C2 => n32, Y => 
                           crossbar_out(154));
   U981 : OAI222xp33_ASAP7_75t_R port map( A1 => n304, A2 => n26, B1 => n240, 
                           B2 => n38, C1 => n930, C2 => n32, Y => 
                           crossbar_out(153));
   U982 : OAI222xp33_ASAP7_75t_R port map( A1 => n305, A2 => n26, B1 => n241, 
                           B2 => n38, C1 => n929, C2 => n32, Y => 
                           crossbar_out(152));
   U983 : OAI222xp33_ASAP7_75t_R port map( A1 => n306, A2 => n26, B1 => n242, 
                           B2 => n38, C1 => n928, C2 => n32, Y => 
                           crossbar_out(151));
   U984 : OAI222xp33_ASAP7_75t_R port map( A1 => n307, A2 => n26, B1 => n243, 
                           B2 => n38, C1 => n927, C2 => n32, Y => 
                           crossbar_out(150));
   U985 : OAI222xp33_ASAP7_75t_R port map( A1 => n308, A2 => n26, B1 => n244, 
                           B2 => n38, C1 => n926, C2 => n32, Y => 
                           crossbar_out(149));
   U986 : OAI222xp33_ASAP7_75t_R port map( A1 => n309, A2 => n26, B1 => n245, 
                           B2 => n38, C1 => n925, C2 => n32, Y => 
                           crossbar_out(148));
   U987 : OAI222xp33_ASAP7_75t_R port map( A1 => n328, A2 => n25, B1 => n264, 
                           B2 => n37, C1 => n924, C2 => n31, Y => 
                           crossbar_out(129));
   U988 : OAI222xp33_ASAP7_75t_R port map( A1 => n310, A2 => n25, B1 => n246, 
                           B2 => n37, C1 => n923, C2 => n31, Y => 
                           crossbar_out(147));
   U989 : OAI222xp33_ASAP7_75t_R port map( A1 => n311, A2 => n25, B1 => n247, 
                           B2 => n37, C1 => n922, C2 => n31, Y => 
                           crossbar_out(146));
   U990 : OAI222xp33_ASAP7_75t_R port map( A1 => n312, A2 => n25, B1 => n248, 
                           B2 => n37, C1 => n921, C2 => n31, Y => 
                           crossbar_out(145));
   U991 : OAI222xp33_ASAP7_75t_R port map( A1 => n313, A2 => n25, B1 => n249, 
                           B2 => n37, C1 => n920, C2 => n31, Y => 
                           crossbar_out(144));
   U992 : OAI222xp33_ASAP7_75t_R port map( A1 => n314, A2 => n25, B1 => n250, 
                           B2 => n37, C1 => n919, C2 => n31, Y => 
                           crossbar_out(143));
   U993 : OAI222xp33_ASAP7_75t_R port map( A1 => n315, A2 => n25, B1 => n251, 
                           B2 => n37, C1 => n918, C2 => n31, Y => 
                           crossbar_out(142));
   U994 : OAI222xp33_ASAP7_75t_R port map( A1 => n316, A2 => n25, B1 => n252, 
                           B2 => n37, C1 => n917, C2 => n31, Y => 
                           crossbar_out(141));
   U995 : OAI222xp33_ASAP7_75t_R port map( A1 => n317, A2 => n25, B1 => n253, 
                           B2 => n37, C1 => n916, C2 => n31, Y => 
                           crossbar_out(140));
   U996 : OAI222xp33_ASAP7_75t_R port map( A1 => n318, A2 => n25, B1 => n254, 
                           B2 => n37, C1 => n915, C2 => n31, Y => 
                           crossbar_out(139));
   U997 : OAI222xp33_ASAP7_75t_R port map( A1 => n319, A2 => n25, B1 => n255, 
                           B2 => n37, C1 => n914, C2 => n31, Y => 
                           crossbar_out(138));
   U998 : OAI222xp33_ASAP7_75t_R port map( A1 => n329, A2 => n25, B1 => n265, 
                           B2 => n37, C1 => n913, C2 => n31, Y => 
                           crossbar_out(128));
   U999 : OAI221xp5_ASAP7_75t_R port map( A1 => n853, A2 => n96, B1 => n976, B2
                           => n24, C => n607, Y => crossbar_out(73));
   U1000 : AOI222xp33_ASAP7_75t_R port map( A1 => n90, A2 => crossbar_in(201), 
                           B1 => n84, B2 => crossbar_in(329), C1 => n78, C2 => 
                           crossbar_in(265), Y => n607);
   U1001 : OAI221xp5_ASAP7_75t_R port map( A1 => n854, A2 => n96, B1 => n975, 
                           B2 => n24, C => n611, Y => crossbar_out(72));
   U1002 : AOI222xp33_ASAP7_75t_R port map( A1 => n90, A2 => crossbar_in(200), 
                           B1 => n84, B2 => crossbar_in(328), C1 => n78, C2 => 
                           crossbar_in(264), Y => n611);
   U1003 : OAI221xp5_ASAP7_75t_R port map( A1 => n855, A2 => n96, B1 => n974, 
                           B2 => n24, C => n612, Y => crossbar_out(71));
   U1004 : AOI222xp33_ASAP7_75t_R port map( A1 => n90, A2 => crossbar_in(199), 
                           B1 => n84, B2 => crossbar_in(327), C1 => n78, C2 => 
                           crossbar_in(263), Y => n612);
   U1005 : OAI221xp5_ASAP7_75t_R port map( A1 => n856, A2 => n96, B1 => n973, 
                           B2 => n24, C => n613, Y => crossbar_out(70));
   U1006 : AOI222xp33_ASAP7_75t_R port map( A1 => n90, A2 => crossbar_in(198), 
                           B1 => n84, B2 => crossbar_in(326), C1 => n78, C2 => 
                           crossbar_in(262), Y => n613);
   U1007 : OAI221xp5_ASAP7_75t_R port map( A1 => n863, A2 => n96, B1 => n972, 
                           B2 => n23, C => n614, Y => crossbar_out(127));
   U1008 : AOI222xp33_ASAP7_75t_R port map( A1 => n90, A2 => crossbar_in(255), 
                           B1 => n84, B2 => crossbar_in(383), C1 => n78, C2 => 
                           crossbar_in(319), Y => n614);
   U1009 : OAI221xp5_ASAP7_75t_R port map( A1 => n864, A2 => n96, B1 => n971, 
                           B2 => n23, C => n615, Y => crossbar_out(126));
   U1010 : AOI222xp33_ASAP7_75t_R port map( A1 => n90, A2 => crossbar_in(254), 
                           B1 => n84, B2 => crossbar_in(382), C1 => n78, C2 => 
                           crossbar_in(318), Y => n615);
   U1011 : OAI221xp5_ASAP7_75t_R port map( A1 => n865, A2 => n96, B1 => n970, 
                           B2 => n23, C => n616, Y => crossbar_out(125));
   U1012 : AOI222xp33_ASAP7_75t_R port map( A1 => n90, A2 => crossbar_in(253), 
                           B1 => n84, B2 => crossbar_in(381), C1 => n78, C2 => 
                           crossbar_in(317), Y => n616);
   U1013 : OAI221xp5_ASAP7_75t_R port map( A1 => n866, A2 => n96, B1 => n969, 
                           B2 => n23, C => n617, Y => crossbar_out(124));
   U1014 : AOI222xp33_ASAP7_75t_R port map( A1 => n90, A2 => crossbar_in(252), 
                           B1 => n84, B2 => crossbar_in(380), C1 => n78, C2 => 
                           crossbar_in(316), Y => n617);
   U1015 : OAI221xp5_ASAP7_75t_R port map( A1 => n857, A2 => n96, B1 => n968, 
                           B2 => n23, C => n618, Y => crossbar_out(69));
   U1016 : AOI222xp33_ASAP7_75t_R port map( A1 => n90, A2 => crossbar_in(197), 
                           B1 => n84, B2 => crossbar_in(325), C1 => n78, C2 => 
                           crossbar_in(261), Y => n618);
   U1017 : OAI221xp5_ASAP7_75t_R port map( A1 => n867, A2 => n96, B1 => n967, 
                           B2 => n23, C => n619, Y => crossbar_out(123));
   U1018 : AOI222xp33_ASAP7_75t_R port map( A1 => n90, A2 => crossbar_in(251), 
                           B1 => n84, B2 => crossbar_in(379), C1 => n78, C2 => 
                           crossbar_in(315), Y => n619);
   U1019 : OAI221xp5_ASAP7_75t_R port map( A1 => n868, A2 => n96, B1 => n966, 
                           B2 => n23, C => n620, Y => crossbar_out(122));
   U1020 : AOI222xp33_ASAP7_75t_R port map( A1 => n90, A2 => crossbar_in(250), 
                           B1 => n84, B2 => crossbar_in(378), C1 => n78, C2 => 
                           crossbar_in(314), Y => n620);
   U1021 : OAI221xp5_ASAP7_75t_R port map( A1 => n869, A2 => n96, B1 => n965, 
                           B2 => n23, C => n621, Y => crossbar_out(121));
   U1022 : AOI222xp33_ASAP7_75t_R port map( A1 => n90, A2 => crossbar_in(249), 
                           B1 => n84, B2 => crossbar_in(377), C1 => n78, C2 => 
                           crossbar_in(313), Y => n621);
   U1023 : OAI221xp5_ASAP7_75t_R port map( A1 => n870, A2 => n97, B1 => n964, 
                           B2 => n23, C => n622, Y => crossbar_out(120));
   U1024 : AOI222xp33_ASAP7_75t_R port map( A1 => n91, A2 => crossbar_in(248), 
                           B1 => n85, B2 => crossbar_in(376), C1 => n79, C2 => 
                           crossbar_in(312), Y => n622);
   U1025 : OAI221xp5_ASAP7_75t_R port map( A1 => n871, A2 => n97, B1 => n963, 
                           B2 => n23, C => n623, Y => crossbar_out(119));
   U1026 : AOI222xp33_ASAP7_75t_R port map( A1 => n91, A2 => crossbar_in(247), 
                           B1 => n85, B2 => crossbar_in(375), C1 => n79, C2 => 
                           crossbar_in(311), Y => n623);
   U1027 : OAI221xp5_ASAP7_75t_R port map( A1 => n872, A2 => n97, B1 => n962, 
                           B2 => n23, C => n624, Y => crossbar_out(118));
   U1028 : AOI222xp33_ASAP7_75t_R port map( A1 => n91, A2 => crossbar_in(246), 
                           B1 => n85, B2 => crossbar_in(374), C1 => n79, C2 => 
                           crossbar_in(310), Y => n624);
   U1029 : OAI221xp5_ASAP7_75t_R port map( A1 => n873, A2 => n97, B1 => n961, 
                           B2 => n23, C => n625, Y => crossbar_out(117));
   U1030 : AOI222xp33_ASAP7_75t_R port map( A1 => n91, A2 => crossbar_in(245), 
                           B1 => n85, B2 => crossbar_in(373), C1 => n79, C2 => 
                           crossbar_in(309), Y => n625);
   U1031 : OAI221xp5_ASAP7_75t_R port map( A1 => n874, A2 => n97, B1 => n960, 
                           B2 => n22, C => n626, Y => crossbar_out(116));
   U1032 : AOI222xp33_ASAP7_75t_R port map( A1 => n91, A2 => crossbar_in(244), 
                           B1 => n85, B2 => crossbar_in(372), C1 => n79, C2 => 
                           crossbar_in(308), Y => n626);
   U1033 : OAI221xp5_ASAP7_75t_R port map( A1 => n875, A2 => n97, B1 => n959, 
                           B2 => n22, C => n627, Y => crossbar_out(115));
   U1034 : AOI222xp33_ASAP7_75t_R port map( A1 => n91, A2 => crossbar_in(243), 
                           B1 => n85, B2 => crossbar_in(371), C1 => n79, C2 => 
                           crossbar_in(307), Y => n627);
   U1035 : OAI221xp5_ASAP7_75t_R port map( A1 => n876, A2 => n97, B1 => n958, 
                           B2 => n22, C => n628, Y => crossbar_out(114));
   U1036 : AOI222xp33_ASAP7_75t_R port map( A1 => n91, A2 => crossbar_in(242), 
                           B1 => n85, B2 => crossbar_in(370), C1 => n79, C2 => 
                           crossbar_in(306), Y => n628);
   U1037 : OAI221xp5_ASAP7_75t_R port map( A1 => n858, A2 => n97, B1 => n957, 
                           B2 => n22, C => n629, Y => crossbar_out(68));
   U1038 : AOI222xp33_ASAP7_75t_R port map( A1 => n91, A2 => crossbar_in(196), 
                           B1 => n85, B2 => crossbar_in(324), C1 => n79, C2 => 
                           crossbar_in(260), Y => n629);
   U1039 : OAI221xp5_ASAP7_75t_R port map( A1 => n877, A2 => n97, B1 => n956, 
                           B2 => n22, C => n630, Y => crossbar_out(113));
   U1040 : AOI222xp33_ASAP7_75t_R port map( A1 => n91, A2 => crossbar_in(241), 
                           B1 => n85, B2 => crossbar_in(369), C1 => n79, C2 => 
                           crossbar_in(305), Y => n630);
   U1041 : OAI221xp5_ASAP7_75t_R port map( A1 => n878, A2 => n97, B1 => n955, 
                           B2 => n22, C => n631, Y => crossbar_out(112));
   U1042 : AOI222xp33_ASAP7_75t_R port map( A1 => n91, A2 => crossbar_in(240), 
                           B1 => n85, B2 => crossbar_in(368), C1 => n79, C2 => 
                           crossbar_in(304), Y => n631);
   U1043 : OAI221xp5_ASAP7_75t_R port map( A1 => n879, A2 => n97, B1 => n954, 
                           B2 => n22, C => n632, Y => crossbar_out(111));
   U1044 : AOI222xp33_ASAP7_75t_R port map( A1 => n91, A2 => crossbar_in(239), 
                           B1 => n85, B2 => crossbar_in(367), C1 => n79, C2 => 
                           crossbar_in(303), Y => n632);
   U1045 : OAI221xp5_ASAP7_75t_R port map( A1 => n880, A2 => n97, B1 => n953, 
                           B2 => n22, C => n633, Y => crossbar_out(110));
   U1046 : AOI222xp33_ASAP7_75t_R port map( A1 => n91, A2 => crossbar_in(238), 
                           B1 => n85, B2 => crossbar_in(366), C1 => n79, C2 => 
                           crossbar_in(302), Y => n633);
   U1047 : OAI221xp5_ASAP7_75t_R port map( A1 => n881, A2 => n98, B1 => n952, 
                           B2 => n22, C => n634, Y => crossbar_out(109));
   U1048 : AOI222xp33_ASAP7_75t_R port map( A1 => n92, A2 => crossbar_in(237), 
                           B1 => n86, B2 => crossbar_in(365), C1 => n80, C2 => 
                           crossbar_in(301), Y => n634);
   U1049 : OAI221xp5_ASAP7_75t_R port map( A1 => n882, A2 => n98, B1 => n951, 
                           B2 => n22, C => n635, Y => crossbar_out(108));
   U1050 : AOI222xp33_ASAP7_75t_R port map( A1 => n92, A2 => crossbar_in(236), 
                           B1 => n86, B2 => crossbar_in(364), C1 => n80, C2 => 
                           crossbar_in(300), Y => n635);
   U1051 : OAI221xp5_ASAP7_75t_R port map( A1 => n883, A2 => n98, B1 => n950, 
                           B2 => n22, C => n636, Y => crossbar_out(107));
   U1052 : AOI222xp33_ASAP7_75t_R port map( A1 => n92, A2 => crossbar_in(235), 
                           B1 => n86, B2 => crossbar_in(363), C1 => n80, C2 => 
                           crossbar_in(299), Y => n636);
   U1053 : OAI221xp5_ASAP7_75t_R port map( A1 => n884, A2 => n98, B1 => n949, 
                           B2 => n22, C => n637, Y => crossbar_out(106));
   U1054 : AOI222xp33_ASAP7_75t_R port map( A1 => n92, A2 => crossbar_in(234), 
                           B1 => n86, B2 => crossbar_in(362), C1 => n80, C2 => 
                           crossbar_in(298), Y => n637);
   U1055 : OAI221xp5_ASAP7_75t_R port map( A1 => n885, A2 => n98, B1 => n948, 
                           B2 => n21, C => n638, Y => crossbar_out(105));
   U1056 : AOI222xp33_ASAP7_75t_R port map( A1 => n92, A2 => crossbar_in(233), 
                           B1 => n86, B2 => crossbar_in(361), C1 => n80, C2 => 
                           crossbar_in(297), Y => n638);
   U1057 : OAI221xp5_ASAP7_75t_R port map( A1 => n886, A2 => n98, B1 => n947, 
                           B2 => n21, C => n639, Y => crossbar_out(104));
   U1058 : AOI222xp33_ASAP7_75t_R port map( A1 => n92, A2 => crossbar_in(232), 
                           B1 => n86, B2 => crossbar_in(360), C1 => n80, C2 => 
                           crossbar_in(296), Y => n639);
   U1059 : OAI221xp5_ASAP7_75t_R port map( A1 => n859, A2 => n98, B1 => n946, 
                           B2 => n21, C => n640, Y => crossbar_out(67));
   U1060 : AOI222xp33_ASAP7_75t_R port map( A1 => n92, A2 => crossbar_in(195), 
                           B1 => n86, B2 => crossbar_in(323), C1 => n80, C2 => 
                           crossbar_in(259), Y => n640);
   U1061 : OAI221xp5_ASAP7_75t_R port map( A1 => n887, A2 => n98, B1 => n945, 
                           B2 => n21, C => n641, Y => crossbar_out(103));
   U1062 : AOI222xp33_ASAP7_75t_R port map( A1 => n92, A2 => crossbar_in(231), 
                           B1 => n86, B2 => crossbar_in(359), C1 => n80, C2 => 
                           crossbar_in(295), Y => n641);
   U1063 : OAI221xp5_ASAP7_75t_R port map( A1 => n888, A2 => n98, B1 => n944, 
                           B2 => n21, C => n642, Y => crossbar_out(102));
   U1064 : AOI222xp33_ASAP7_75t_R port map( A1 => n92, A2 => crossbar_in(230), 
                           B1 => n86, B2 => crossbar_in(358), C1 => n80, C2 => 
                           crossbar_in(294), Y => n642);
   U1065 : OAI221xp5_ASAP7_75t_R port map( A1 => n889, A2 => n98, B1 => n943, 
                           B2 => n21, C => n643, Y => crossbar_out(101));
   U1066 : AOI222xp33_ASAP7_75t_R port map( A1 => n92, A2 => crossbar_in(229), 
                           B1 => n86, B2 => crossbar_in(357), C1 => n80, C2 => 
                           crossbar_in(293), Y => n643);
   U1067 : OAI221xp5_ASAP7_75t_R port map( A1 => n890, A2 => n98, B1 => n942, 
                           B2 => n21, C => n644, Y => crossbar_out(100));
   U1068 : AOI222xp33_ASAP7_75t_R port map( A1 => n92, A2 => crossbar_in(228), 
                           B1 => n86, B2 => crossbar_in(356), C1 => n80, C2 => 
                           crossbar_in(292), Y => n644);
   U1069 : OAI221xp5_ASAP7_75t_R port map( A1 => n891, A2 => n98, B1 => n941, 
                           B2 => n21, C => n645, Y => crossbar_out(99));
   U1070 : AOI222xp33_ASAP7_75t_R port map( A1 => n92, A2 => crossbar_in(227), 
                           B1 => n86, B2 => crossbar_in(355), C1 => n80, C2 => 
                           crossbar_in(291), Y => n645);
   U1071 : OAI221xp5_ASAP7_75t_R port map( A1 => n892, A2 => n99, B1 => n940, 
                           B2 => n21, C => n646, Y => crossbar_out(98));
   U1072 : AOI222xp33_ASAP7_75t_R port map( A1 => n93, A2 => crossbar_in(226), 
                           B1 => n87, B2 => crossbar_in(354), C1 => n81, C2 => 
                           crossbar_in(290), Y => n646);
   U1073 : OAI221xp5_ASAP7_75t_R port map( A1 => n893, A2 => n99, B1 => n939, 
                           B2 => n21, C => n647, Y => crossbar_out(97));
   U1074 : AOI222xp33_ASAP7_75t_R port map( A1 => n93, A2 => crossbar_in(225), 
                           B1 => n87, B2 => crossbar_in(353), C1 => n81, C2 => 
                           crossbar_in(289), Y => n647);
   U1075 : OAI221xp5_ASAP7_75t_R port map( A1 => n894, A2 => n99, B1 => n938, 
                           B2 => n21, C => n648, Y => crossbar_out(96));
   U1076 : AOI222xp33_ASAP7_75t_R port map( A1 => n93, A2 => crossbar_in(224), 
                           B1 => n87, B2 => crossbar_in(352), C1 => n81, C2 => 
                           crossbar_in(288), Y => n648);
   U1077 : OAI221xp5_ASAP7_75t_R port map( A1 => n895, A2 => n99, B1 => n937, 
                           B2 => n21, C => n649, Y => crossbar_out(95));
   U1078 : AOI222xp33_ASAP7_75t_R port map( A1 => n93, A2 => crossbar_in(223), 
                           B1 => n87, B2 => crossbar_in(351), C1 => n81, C2 => 
                           crossbar_in(287), Y => n649);
   U1079 : OAI221xp5_ASAP7_75t_R port map( A1 => n896, A2 => n99, B1 => n936, 
                           B2 => n20, C => n650, Y => crossbar_out(94));
   U1080 : AOI222xp33_ASAP7_75t_R port map( A1 => n93, A2 => crossbar_in(222), 
                           B1 => n87, B2 => crossbar_in(350), C1 => n81, C2 => 
                           crossbar_in(286), Y => n650);
   U1081 : OAI221xp5_ASAP7_75t_R port map( A1 => n860, A2 => n99, B1 => n935, 
                           B2 => n20, C => n651, Y => crossbar_out(66));
   U1082 : AOI222xp33_ASAP7_75t_R port map( A1 => n93, A2 => crossbar_in(194), 
                           B1 => n87, B2 => crossbar_in(322), C1 => n81, C2 => 
                           crossbar_in(258), Y => n651);
   U1083 : OAI221xp5_ASAP7_75t_R port map( A1 => n833, A2 => n99, B1 => n934, 
                           B2 => n20, C => n652, Y => crossbar_out(93));
   U1084 : AOI222xp33_ASAP7_75t_R port map( A1 => n93, A2 => crossbar_in(221), 
                           B1 => n87, B2 => crossbar_in(349), C1 => n81, C2 => 
                           crossbar_in(285), Y => n652);
   U1085 : OAI221xp5_ASAP7_75t_R port map( A1 => n834, A2 => n99, B1 => n933, 
                           B2 => n20, C => n653, Y => crossbar_out(92));
   U1086 : AOI222xp33_ASAP7_75t_R port map( A1 => n93, A2 => crossbar_in(220), 
                           B1 => n87, B2 => crossbar_in(348), C1 => n81, C2 => 
                           crossbar_in(284), Y => n653);
   U1087 : OAI221xp5_ASAP7_75t_R port map( A1 => n835, A2 => n99, B1 => n932, 
                           B2 => n20, C => n654, Y => crossbar_out(91));
   U1088 : AOI222xp33_ASAP7_75t_R port map( A1 => n93, A2 => crossbar_in(219), 
                           B1 => n87, B2 => crossbar_in(347), C1 => n81, C2 => 
                           crossbar_in(283), Y => n654);
   U1089 : OAI221xp5_ASAP7_75t_R port map( A1 => n836, A2 => n99, B1 => n931, 
                           B2 => n20, C => n655, Y => crossbar_out(90));
   U1090 : AOI222xp33_ASAP7_75t_R port map( A1 => n93, A2 => crossbar_in(218), 
                           B1 => n87, B2 => crossbar_in(346), C1 => n81, C2 => 
                           crossbar_in(282), Y => n655);
   U1091 : OAI221xp5_ASAP7_75t_R port map( A1 => n837, A2 => n99, B1 => n930, 
                           B2 => n20, C => n656, Y => crossbar_out(89));
   U1092 : AOI222xp33_ASAP7_75t_R port map( A1 => n93, A2 => crossbar_in(217), 
                           B1 => n87, B2 => crossbar_in(345), C1 => n81, C2 => 
                           crossbar_in(281), Y => n656);
   U1093 : OAI221xp5_ASAP7_75t_R port map( A1 => n838, A2 => n99, B1 => n929, 
                           B2 => n20, C => n657, Y => crossbar_out(88));
   U1094 : AOI222xp33_ASAP7_75t_R port map( A1 => n93, A2 => crossbar_in(216), 
                           B1 => n87, B2 => crossbar_in(344), C1 => n81, C2 => 
                           crossbar_in(280), Y => n657);
   U1095 : OAI221xp5_ASAP7_75t_R port map( A1 => n839, A2 => n100, B1 => n928, 
                           B2 => n20, C => n658, Y => crossbar_out(87));
   U1096 : AOI222xp33_ASAP7_75t_R port map( A1 => n94, A2 => crossbar_in(215), 
                           B1 => n88, B2 => crossbar_in(343), C1 => n82, C2 => 
                           crossbar_in(279), Y => n658);
   U1097 : OAI221xp5_ASAP7_75t_R port map( A1 => n840, A2 => n100, B1 => n927, 
                           B2 => n20, C => n659, Y => crossbar_out(86));
   U1098 : AOI222xp33_ASAP7_75t_R port map( A1 => n94, A2 => crossbar_in(214), 
                           B1 => n88, B2 => crossbar_in(342), C1 => n82, C2 => 
                           crossbar_in(278), Y => n659);
   U1099 : OAI221xp5_ASAP7_75t_R port map( A1 => n841, A2 => n100, B1 => n926, 
                           B2 => n20, C => n660, Y => crossbar_out(85));
   U1100 : AOI222xp33_ASAP7_75t_R port map( A1 => n94, A2 => crossbar_in(213), 
                           B1 => n88, B2 => crossbar_in(341), C1 => n82, C2 => 
                           crossbar_in(277), Y => n660);
   U1101 : OAI221xp5_ASAP7_75t_R port map( A1 => n842, A2 => n100, B1 => n925, 
                           B2 => n20, C => n661, Y => crossbar_out(84));
   U1102 : AOI222xp33_ASAP7_75t_R port map( A1 => n94, A2 => crossbar_in(212), 
                           B1 => n88, B2 => crossbar_in(340), C1 => n82, C2 => 
                           crossbar_in(276), Y => n661);
   U1103 : OAI221xp5_ASAP7_75t_R port map( A1 => n861, A2 => n100, B1 => n924, 
                           B2 => n19, C => n662, Y => crossbar_out(65));
   U1104 : AOI222xp33_ASAP7_75t_R port map( A1 => n94, A2 => crossbar_in(193), 
                           B1 => n88, B2 => crossbar_in(321), C1 => n82, C2 => 
                           crossbar_in(257), Y => n662);
   U1105 : OAI221xp5_ASAP7_75t_R port map( A1 => n843, A2 => n100, B1 => n923, 
                           B2 => n19, C => n663, Y => crossbar_out(83));
   U1106 : AOI222xp33_ASAP7_75t_R port map( A1 => n94, A2 => crossbar_in(211), 
                           B1 => n88, B2 => crossbar_in(339), C1 => n82, C2 => 
                           crossbar_in(275), Y => n663);
   U1107 : OAI221xp5_ASAP7_75t_R port map( A1 => n844, A2 => n100, B1 => n922, 
                           B2 => n19, C => n664, Y => crossbar_out(82));
   U1108 : AOI222xp33_ASAP7_75t_R port map( A1 => n94, A2 => crossbar_in(210), 
                           B1 => n88, B2 => crossbar_in(338), C1 => n82, C2 => 
                           crossbar_in(274), Y => n664);
   U1109 : OAI221xp5_ASAP7_75t_R port map( A1 => n845, A2 => n100, B1 => n921, 
                           B2 => n19, C => n665, Y => crossbar_out(81));
   U1110 : AOI222xp33_ASAP7_75t_R port map( A1 => n94, A2 => crossbar_in(209), 
                           B1 => n88, B2 => crossbar_in(337), C1 => n82, C2 => 
                           crossbar_in(273), Y => n665);
   U1111 : OAI221xp5_ASAP7_75t_R port map( A1 => n846, A2 => n100, B1 => n920, 
                           B2 => n19, C => n666, Y => crossbar_out(80));
   U1112 : AOI222xp33_ASAP7_75t_R port map( A1 => n94, A2 => crossbar_in(208), 
                           B1 => n88, B2 => crossbar_in(336), C1 => n82, C2 => 
                           crossbar_in(272), Y => n666);
   U1113 : OAI221xp5_ASAP7_75t_R port map( A1 => n847, A2 => n100, B1 => n919, 
                           B2 => n19, C => n667, Y => crossbar_out(79));
   U1114 : AOI222xp33_ASAP7_75t_R port map( A1 => n94, A2 => crossbar_in(207), 
                           B1 => n88, B2 => crossbar_in(335), C1 => n82, C2 => 
                           crossbar_in(271), Y => n667);
   U1115 : OAI221xp5_ASAP7_75t_R port map( A1 => n848, A2 => n100, B1 => n918, 
                           B2 => n19, C => n668, Y => crossbar_out(78));
   U1116 : AOI222xp33_ASAP7_75t_R port map( A1 => n94, A2 => crossbar_in(206), 
                           B1 => n88, B2 => crossbar_in(334), C1 => n82, C2 => 
                           crossbar_in(270), Y => n668);
   U1117 : OAI221xp5_ASAP7_75t_R port map( A1 => n849, A2 => n100, B1 => n917, 
                           B2 => n19, C => n669, Y => crossbar_out(77));
   U1118 : AOI222xp33_ASAP7_75t_R port map( A1 => n94, A2 => crossbar_in(205), 
                           B1 => n88, B2 => crossbar_in(333), C1 => n82, C2 => 
                           crossbar_in(269), Y => n669);
   U1119 : OAI221xp5_ASAP7_75t_R port map( A1 => n850, A2 => n101, B1 => n916, 
                           B2 => n19, C => n670, Y => crossbar_out(76));
   U1120 : AOI222xp33_ASAP7_75t_R port map( A1 => n95, A2 => crossbar_in(204), 
                           B1 => n89, B2 => crossbar_in(332), C1 => n83, C2 => 
                           crossbar_in(268), Y => n670);
   U1121 : OAI221xp5_ASAP7_75t_R port map( A1 => n851, A2 => n101, B1 => n915, 
                           B2 => n19, C => n671, Y => crossbar_out(75));
   U1122 : AOI222xp33_ASAP7_75t_R port map( A1 => n95, A2 => crossbar_in(203), 
                           B1 => n89, B2 => crossbar_in(331), C1 => n83, C2 => 
                           crossbar_in(267), Y => n671);
   U1123 : OAI221xp5_ASAP7_75t_R port map( A1 => n852, A2 => n101, B1 => n914, 
                           B2 => n19, C => n672, Y => crossbar_out(74));
   U1124 : AOI222xp33_ASAP7_75t_R port map( A1 => n95, A2 => crossbar_in(202), 
                           B1 => n89, B2 => crossbar_in(330), C1 => n83, C2 => 
                           crossbar_in(266), Y => n672);
   U1125 : OAI221xp5_ASAP7_75t_R port map( A1 => n862, A2 => n101, B1 => n913, 
                           B2 => n19, C => n673, Y => crossbar_out(64));
   U1126 : AOI222xp33_ASAP7_75t_R port map( A1 => n95, A2 => crossbar_in(192), 
                           B1 => n89, B2 => crossbar_in(320), C1 => n83, C2 => 
                           crossbar_in(256), Y => n673);
   U1127 : OAI211xp5_ASAP7_75t_R port map( A1 => n192, A2 => n77, B => n675, C 
                           => n676, Y => crossbar_out(9));
   U1128 : AOI222xp33_ASAP7_75t_R port map( A1 => n67, A2 => crossbar_in(265), 
                           B1 => n61, B2 => crossbar_in(393), C1 => n55, C2 => 
                           crossbar_in(329), Y => n676);
   U1129 : OAI211xp5_ASAP7_75t_R port map( A1 => n193, A2 => n77, B => n682, C 
                           => n683, Y => crossbar_out(8));
   U1130 : AOI222xp33_ASAP7_75t_R port map( A1 => n67, A2 => crossbar_in(264), 
                           B1 => n61, B2 => crossbar_in(392), C1 => n55, C2 => 
                           crossbar_in(328), Y => n683);
   U1131 : OAI211xp5_ASAP7_75t_R port map( A1 => n194, A2 => n77, B => n684, C 
                           => n685, Y => crossbar_out(7));
   U1132 : AOI222xp33_ASAP7_75t_R port map( A1 => n67, A2 => crossbar_in(263), 
                           B1 => n61, B2 => crossbar_in(391), C1 => n55, C2 => 
                           crossbar_in(327), Y => n685);
   U1133 : OAI211xp5_ASAP7_75t_R port map( A1 => n195, A2 => n77, B => n686, C 
                           => n687, Y => crossbar_out(6));
   U1134 : AOI222xp33_ASAP7_75t_R port map( A1 => n67, A2 => crossbar_in(262), 
                           B1 => n61, B2 => crossbar_in(390), C1 => n55, C2 => 
                           crossbar_in(326), Y => n687);
   U1135 : OAI211xp5_ASAP7_75t_R port map( A1 => n202, A2 => n77, B => n688, C 
                           => n689, Y => crossbar_out(63));
   U1136 : AOI222xp33_ASAP7_75t_R port map( A1 => n67, A2 => crossbar_in(319), 
                           B1 => n61, B2 => crossbar_in(447), C1 => n55, C2 => 
                           crossbar_in(383), Y => n689);
   U1137 : OAI211xp5_ASAP7_75t_R port map( A1 => n203, A2 => n77, B => n690, C 
                           => n691, Y => crossbar_out(62));
   U1138 : AOI222xp33_ASAP7_75t_R port map( A1 => n67, A2 => crossbar_in(318), 
                           B1 => n61, B2 => crossbar_in(446), C1 => n55, C2 => 
                           crossbar_in(382), Y => n691);
   U1139 : OAI211xp5_ASAP7_75t_R port map( A1 => n204, A2 => n77, B => n692, C 
                           => n693, Y => crossbar_out(61));
   U1140 : AOI222xp33_ASAP7_75t_R port map( A1 => n67, A2 => crossbar_in(317), 
                           B1 => n61, B2 => crossbar_in(445), C1 => n55, C2 => 
                           crossbar_in(381), Y => n693);
   U1141 : OAI211xp5_ASAP7_75t_R port map( A1 => n205, A2 => n77, B => n694, C 
                           => n695, Y => crossbar_out(60));
   U1142 : AOI222xp33_ASAP7_75t_R port map( A1 => n67, A2 => crossbar_in(316), 
                           B1 => n61, B2 => crossbar_in(444), C1 => n55, C2 => 
                           crossbar_in(380), Y => n695);
   U1143 : OAI211xp5_ASAP7_75t_R port map( A1 => n196, A2 => n77, B => n696, C 
                           => n697, Y => crossbar_out(5));
   U1144 : AOI222xp33_ASAP7_75t_R port map( A1 => n67, A2 => crossbar_in(261), 
                           B1 => n61, B2 => crossbar_in(389), C1 => n55, C2 => 
                           crossbar_in(325), Y => n697);
   U1145 : OAI211xp5_ASAP7_75t_R port map( A1 => n206, A2 => n77, B => n698, C 
                           => n699, Y => crossbar_out(59));
   U1146 : AOI222xp33_ASAP7_75t_R port map( A1 => n67, A2 => crossbar_in(315), 
                           B1 => n61, B2 => crossbar_in(443), C1 => n55, C2 => 
                           crossbar_in(379), Y => n699);
   U1147 : OAI211xp5_ASAP7_75t_R port map( A1 => n207, A2 => n77, B => n700, C 
                           => n701, Y => crossbar_out(58));
   U1148 : AOI222xp33_ASAP7_75t_R port map( A1 => n67, A2 => crossbar_in(314), 
                           B1 => n61, B2 => crossbar_in(442), C1 => n55, C2 => 
                           crossbar_in(378), Y => n701);
   U1149 : OAI211xp5_ASAP7_75t_R port map( A1 => n208, A2 => n77, B => n702, C 
                           => n703, Y => crossbar_out(57));
   U1150 : AOI222xp33_ASAP7_75t_R port map( A1 => n67, A2 => crossbar_in(313), 
                           B1 => n61, B2 => crossbar_in(441), C1 => n55, C2 => 
                           crossbar_in(377), Y => n703);
   U1151 : OAI211xp5_ASAP7_75t_R port map( A1 => n209, A2 => n76, B => n704, C 
                           => n705, Y => crossbar_out(56));
   U1152 : AOI222xp33_ASAP7_75t_R port map( A1 => n68, A2 => crossbar_in(312), 
                           B1 => n62, B2 => crossbar_in(440), C1 => n56, C2 => 
                           crossbar_in(376), Y => n705);
   U1153 : OAI211xp5_ASAP7_75t_R port map( A1 => n210, A2 => n76, B => n706, C 
                           => n707, Y => crossbar_out(55));
   U1154 : AOI222xp33_ASAP7_75t_R port map( A1 => n68, A2 => crossbar_in(311), 
                           B1 => n62, B2 => crossbar_in(439), C1 => n56, C2 => 
                           crossbar_in(375), Y => n707);
   U1155 : OAI211xp5_ASAP7_75t_R port map( A1 => n211, A2 => n76, B => n708, C 
                           => n709, Y => crossbar_out(54));
   U1156 : AOI222xp33_ASAP7_75t_R port map( A1 => n68, A2 => crossbar_in(310), 
                           B1 => n62, B2 => crossbar_in(438), C1 => n56, C2 => 
                           crossbar_in(374), Y => n709);
   U1157 : OAI211xp5_ASAP7_75t_R port map( A1 => n212, A2 => n76, B => n710, C 
                           => n711, Y => crossbar_out(53));
   U1158 : AOI222xp33_ASAP7_75t_R port map( A1 => n68, A2 => crossbar_in(309), 
                           B1 => n62, B2 => crossbar_in(437), C1 => n56, C2 => 
                           crossbar_in(373), Y => n711);
   U1159 : OAI211xp5_ASAP7_75t_R port map( A1 => n213, A2 => n76, B => n712, C 
                           => n713, Y => crossbar_out(52));
   U1160 : AOI222xp33_ASAP7_75t_R port map( A1 => n68, A2 => crossbar_in(308), 
                           B1 => n62, B2 => crossbar_in(436), C1 => n56, C2 => 
                           crossbar_in(372), Y => n713);
   U1161 : OAI211xp5_ASAP7_75t_R port map( A1 => n214, A2 => n76, B => n714, C 
                           => n715, Y => crossbar_out(51));
   U1162 : AOI222xp33_ASAP7_75t_R port map( A1 => n68, A2 => crossbar_in(307), 
                           B1 => n62, B2 => crossbar_in(435), C1 => n56, C2 => 
                           crossbar_in(371), Y => n715);
   U1163 : OAI211xp5_ASAP7_75t_R port map( A1 => n215, A2 => n76, B => n716, C 
                           => n717, Y => crossbar_out(50));
   U1164 : AOI222xp33_ASAP7_75t_R port map( A1 => n68, A2 => crossbar_in(306), 
                           B1 => n62, B2 => crossbar_in(434), C1 => n56, C2 => 
                           crossbar_in(370), Y => n717);
   U1165 : OAI211xp5_ASAP7_75t_R port map( A1 => n197, A2 => n76, B => n718, C 
                           => n719, Y => crossbar_out(4));
   U1166 : AOI222xp33_ASAP7_75t_R port map( A1 => n68, A2 => crossbar_in(260), 
                           B1 => n62, B2 => crossbar_in(388), C1 => n56, C2 => 
                           crossbar_in(324), Y => n719);
   U1167 : OAI211xp5_ASAP7_75t_R port map( A1 => n216, A2 => n76, B => n720, C 
                           => n721, Y => crossbar_out(49));
   U1168 : AOI222xp33_ASAP7_75t_R port map( A1 => n68, A2 => crossbar_in(305), 
                           B1 => n62, B2 => crossbar_in(433), C1 => n56, C2 => 
                           crossbar_in(369), Y => n721);
   U1169 : OAI211xp5_ASAP7_75t_R port map( A1 => n217, A2 => n76, B => n722, C 
                           => n723, Y => crossbar_out(48));
   U1170 : AOI222xp33_ASAP7_75t_R port map( A1 => n68, A2 => crossbar_in(304), 
                           B1 => n62, B2 => crossbar_in(432), C1 => n56, C2 => 
                           crossbar_in(368), Y => n723);
   U1171 : OAI211xp5_ASAP7_75t_R port map( A1 => n218, A2 => n76, B => n724, C 
                           => n725, Y => crossbar_out(47));
   U1172 : AOI222xp33_ASAP7_75t_R port map( A1 => n68, A2 => crossbar_in(303), 
                           B1 => n62, B2 => crossbar_in(431), C1 => n56, C2 => 
                           crossbar_in(367), Y => n725);
   U1173 : OAI211xp5_ASAP7_75t_R port map( A1 => n219, A2 => n76, B => n726, C 
                           => n727, Y => crossbar_out(46));
   U1174 : AOI222xp33_ASAP7_75t_R port map( A1 => n68, A2 => crossbar_in(302), 
                           B1 => n62, B2 => crossbar_in(430), C1 => n56, C2 => 
                           crossbar_in(366), Y => n727);
   U1175 : OAI211xp5_ASAP7_75t_R port map( A1 => n220, A2 => n76, B => n728, C 
                           => n729, Y => crossbar_out(45));
   U1176 : AOI222xp33_ASAP7_75t_R port map( A1 => n69, A2 => crossbar_in(301), 
                           B1 => n63, B2 => crossbar_in(429), C1 => n57, C2 => 
                           crossbar_in(365), Y => n729);
   U1177 : OAI211xp5_ASAP7_75t_R port map( A1 => n221, A2 => n75, B => n730, C 
                           => n731, Y => crossbar_out(44));
   U1178 : AOI222xp33_ASAP7_75t_R port map( A1 => n69, A2 => crossbar_in(300), 
                           B1 => n63, B2 => crossbar_in(428), C1 => n57, C2 => 
                           crossbar_in(364), Y => n731);
   U1179 : OAI211xp5_ASAP7_75t_R port map( A1 => n222, A2 => n75, B => n732, C 
                           => n733, Y => crossbar_out(43));
   U1180 : AOI222xp33_ASAP7_75t_R port map( A1 => n69, A2 => crossbar_in(299), 
                           B1 => n63, B2 => crossbar_in(427), C1 => n57, C2 => 
                           crossbar_in(363), Y => n733);
   U1181 : OAI211xp5_ASAP7_75t_R port map( A1 => n223, A2 => n75, B => n734, C 
                           => n735, Y => crossbar_out(42));
   U1182 : AOI222xp33_ASAP7_75t_R port map( A1 => n69, A2 => crossbar_in(298), 
                           B1 => n63, B2 => crossbar_in(426), C1 => n57, C2 => 
                           crossbar_in(362), Y => n735);
   U1183 : OAI211xp5_ASAP7_75t_R port map( A1 => n224, A2 => n75, B => n736, C 
                           => n737, Y => crossbar_out(41));
   U1184 : AOI222xp33_ASAP7_75t_R port map( A1 => n69, A2 => crossbar_in(297), 
                           B1 => n63, B2 => crossbar_in(425), C1 => n57, C2 => 
                           crossbar_in(361), Y => n737);
   U1185 : OAI211xp5_ASAP7_75t_R port map( A1 => n225, A2 => n75, B => n738, C 
                           => n739, Y => crossbar_out(40));
   U1186 : AOI222xp33_ASAP7_75t_R port map( A1 => n69, A2 => crossbar_in(296), 
                           B1 => n63, B2 => crossbar_in(424), C1 => n57, C2 => 
                           crossbar_in(360), Y => n739);
   U1187 : OAI211xp5_ASAP7_75t_R port map( A1 => n198, A2 => n75, B => n740, C 
                           => n741, Y => crossbar_out(3));
   U1188 : AOI222xp33_ASAP7_75t_R port map( A1 => n69, A2 => crossbar_in(259), 
                           B1 => n63, B2 => crossbar_in(387), C1 => n57, C2 => 
                           crossbar_in(323), Y => n741);
   U1189 : OAI211xp5_ASAP7_75t_R port map( A1 => n226, A2 => n75, B => n742, C 
                           => n743, Y => crossbar_out(39));
   U1190 : AOI222xp33_ASAP7_75t_R port map( A1 => n69, A2 => crossbar_in(295), 
                           B1 => n63, B2 => crossbar_in(423), C1 => n57, C2 => 
                           crossbar_in(359), Y => n743);
   U1191 : OAI211xp5_ASAP7_75t_R port map( A1 => n227, A2 => n75, B => n744, C 
                           => n745, Y => crossbar_out(38));
   U1192 : AOI222xp33_ASAP7_75t_R port map( A1 => n69, A2 => crossbar_in(294), 
                           B1 => n63, B2 => crossbar_in(422), C1 => n57, C2 => 
                           crossbar_in(358), Y => n745);
   U1193 : OAI211xp5_ASAP7_75t_R port map( A1 => n228, A2 => n75, B => n746, C 
                           => n747, Y => crossbar_out(37));
   U1194 : AOI222xp33_ASAP7_75t_R port map( A1 => n69, A2 => crossbar_in(293), 
                           B1 => n63, B2 => crossbar_in(421), C1 => n57, C2 => 
                           crossbar_in(357), Y => n747);
   U1195 : OAI211xp5_ASAP7_75t_R port map( A1 => n229, A2 => n75, B => n748, C 
                           => n749, Y => crossbar_out(36));
   U1196 : AOI222xp33_ASAP7_75t_R port map( A1 => n69, A2 => crossbar_in(292), 
                           B1 => n63, B2 => crossbar_in(420), C1 => n57, C2 => 
                           crossbar_in(356), Y => n749);
   U1197 : OAI211xp5_ASAP7_75t_R port map( A1 => n230, A2 => n75, B => n750, C 
                           => n751, Y => crossbar_out(35));
   U1198 : AOI222xp33_ASAP7_75t_R port map( A1 => n69, A2 => crossbar_in(291), 
                           B1 => n63, B2 => crossbar_in(419), C1 => n57, C2 => 
                           crossbar_in(355), Y => n751);
   U1199 : OAI211xp5_ASAP7_75t_R port map( A1 => n231, A2 => n75, B => n752, C 
                           => n753, Y => crossbar_out(34));
   U1200 : AOI222xp33_ASAP7_75t_R port map( A1 => n70, A2 => crossbar_in(290), 
                           B1 => n64, B2 => crossbar_in(418), C1 => n58, C2 => 
                           crossbar_in(354), Y => n753);
   U1201 : OAI211xp5_ASAP7_75t_R port map( A1 => n232, A2 => n75, B => n754, C 
                           => n755, Y => crossbar_out(33));
   U1202 : AOI222xp33_ASAP7_75t_R port map( A1 => n70, A2 => crossbar_in(289), 
                           B1 => n64, B2 => crossbar_in(417), C1 => n58, C2 => 
                           crossbar_in(353), Y => n755);
   U1203 : OAI211xp5_ASAP7_75t_R port map( A1 => n233, A2 => n74, B => n756, C 
                           => n757, Y => crossbar_out(32));
   U1204 : AOI222xp33_ASAP7_75t_R port map( A1 => n70, A2 => crossbar_in(288), 
                           B1 => n64, B2 => crossbar_in(416), C1 => n58, C2 => 
                           crossbar_in(352), Y => n757);
   U1205 : OAI211xp5_ASAP7_75t_R port map( A1 => n234, A2 => n74, B => n758, C 
                           => n759, Y => crossbar_out(31));
   U1206 : AOI222xp33_ASAP7_75t_R port map( A1 => n70, A2 => crossbar_in(287), 
                           B1 => n64, B2 => crossbar_in(415), C1 => n58, C2 => 
                           crossbar_in(351), Y => n759);
   U1207 : OAI211xp5_ASAP7_75t_R port map( A1 => n235, A2 => n74, B => n760, C 
                           => n761, Y => crossbar_out(30));
   U1208 : AOI222xp33_ASAP7_75t_R port map( A1 => n70, A2 => crossbar_in(286), 
                           B1 => n64, B2 => crossbar_in(414), C1 => n58, C2 => 
                           crossbar_in(350), Y => n761);
   U1209 : OAI211xp5_ASAP7_75t_R port map( A1 => n199, A2 => n74, B => n762, C 
                           => n763, Y => crossbar_out(2));
   U1210 : AOI222xp33_ASAP7_75t_R port map( A1 => n70, A2 => crossbar_in(258), 
                           B1 => n64, B2 => crossbar_in(386), C1 => n58, C2 => 
                           crossbar_in(322), Y => n763);
   U1211 : OAI211xp5_ASAP7_75t_R port map( A1 => n172, A2 => n74, B => n764, C 
                           => n765, Y => crossbar_out(29));
   U1212 : AOI222xp33_ASAP7_75t_R port map( A1 => n70, A2 => crossbar_in(285), 
                           B1 => n64, B2 => crossbar_in(413), C1 => n58, C2 => 
                           crossbar_in(349), Y => n765);
   U1213 : OAI211xp5_ASAP7_75t_R port map( A1 => n173, A2 => n74, B => n766, C 
                           => n767, Y => crossbar_out(28));
   U1214 : AOI222xp33_ASAP7_75t_R port map( A1 => n70, A2 => crossbar_in(284), 
                           B1 => n64, B2 => crossbar_in(412), C1 => n58, C2 => 
                           crossbar_in(348), Y => n767);
   U1215 : OAI211xp5_ASAP7_75t_R port map( A1 => n174, A2 => n74, B => n768, C 
                           => n769, Y => crossbar_out(27));
   U1216 : AOI222xp33_ASAP7_75t_R port map( A1 => n70, A2 => crossbar_in(283), 
                           B1 => n64, B2 => crossbar_in(411), C1 => n58, C2 => 
                           crossbar_in(347), Y => n769);
   U1217 : OAI211xp5_ASAP7_75t_R port map( A1 => n175, A2 => n74, B => n770, C 
                           => n771, Y => crossbar_out(26));
   U1218 : AOI222xp33_ASAP7_75t_R port map( A1 => n70, A2 => crossbar_in(282), 
                           B1 => n64, B2 => crossbar_in(410), C1 => n58, C2 => 
                           crossbar_in(346), Y => n771);
   U1219 : OAI211xp5_ASAP7_75t_R port map( A1 => n176, A2 => n74, B => n772, C 
                           => n773, Y => crossbar_out(25));
   U1220 : AOI222xp33_ASAP7_75t_R port map( A1 => n70, A2 => crossbar_in(281), 
                           B1 => n64, B2 => crossbar_in(409), C1 => n58, C2 => 
                           crossbar_in(345), Y => n773);
   U1221 : OAI211xp5_ASAP7_75t_R port map( A1 => n177, A2 => n74, B => n774, C 
                           => n775, Y => crossbar_out(24));
   U1222 : AOI222xp33_ASAP7_75t_R port map( A1 => n70, A2 => crossbar_in(280), 
                           B1 => n64, B2 => crossbar_in(408), C1 => n58, C2 => 
                           crossbar_in(344), Y => n775);
   U1223 : OAI211xp5_ASAP7_75t_R port map( A1 => n178, A2 => n74, B => n776, C 
                           => n777, Y => crossbar_out(23));
   U1224 : AOI222xp33_ASAP7_75t_R port map( A1 => n71, A2 => crossbar_in(279), 
                           B1 => n65, B2 => crossbar_in(407), C1 => n59, C2 => 
                           crossbar_in(343), Y => n777);
   U1225 : OAI211xp5_ASAP7_75t_R port map( A1 => n179, A2 => n74, B => n778, C 
                           => n779, Y => crossbar_out(22));
   U1226 : AOI222xp33_ASAP7_75t_R port map( A1 => n71, A2 => crossbar_in(278), 
                           B1 => n65, B2 => crossbar_in(406), C1 => n59, C2 => 
                           crossbar_in(342), Y => n779);
   U1227 : OAI211xp5_ASAP7_75t_R port map( A1 => n180, A2 => n74, B => n780, C 
                           => n781, Y => crossbar_out(21));
   U1228 : AOI222xp33_ASAP7_75t_R port map( A1 => n71, A2 => crossbar_in(277), 
                           B1 => n65, B2 => crossbar_in(405), C1 => n59, C2 => 
                           crossbar_in(341), Y => n781);
   U1229 : OAI211xp5_ASAP7_75t_R port map( A1 => n181, A2 => n73, B => n782, C 
                           => n783, Y => crossbar_out(20));
   U1230 : AOI222xp33_ASAP7_75t_R port map( A1 => n71, A2 => crossbar_in(276), 
                           B1 => n65, B2 => crossbar_in(404), C1 => n59, C2 => 
                           crossbar_in(340), Y => n783);
   U1231 : OAI211xp5_ASAP7_75t_R port map( A1 => n200, A2 => n73, B => n784, C 
                           => n785, Y => crossbar_out(1));
   U1232 : AOI222xp33_ASAP7_75t_R port map( A1 => n71, A2 => crossbar_in(257), 
                           B1 => n65, B2 => crossbar_in(385), C1 => n59, C2 => 
                           crossbar_in(321), Y => n785);
   U1233 : OAI211xp5_ASAP7_75t_R port map( A1 => n182, A2 => n73, B => n786, C 
                           => n787, Y => crossbar_out(19));
   U1234 : AOI222xp33_ASAP7_75t_R port map( A1 => n71, A2 => crossbar_in(275), 
                           B1 => n65, B2 => crossbar_in(403), C1 => n59, C2 => 
                           crossbar_in(339), Y => n787);
   U1235 : OAI211xp5_ASAP7_75t_R port map( A1 => n183, A2 => n73, B => n788, C 
                           => n789, Y => crossbar_out(18));
   U1236 : AOI222xp33_ASAP7_75t_R port map( A1 => n71, A2 => crossbar_in(274), 
                           B1 => n65, B2 => crossbar_in(402), C1 => n59, C2 => 
                           crossbar_in(338), Y => n789);
   U1237 : OAI211xp5_ASAP7_75t_R port map( A1 => n184, A2 => n73, B => n790, C 
                           => n791, Y => crossbar_out(17));
   U1238 : AOI222xp33_ASAP7_75t_R port map( A1 => n71, A2 => crossbar_in(273), 
                           B1 => n65, B2 => crossbar_in(401), C1 => n59, C2 => 
                           crossbar_in(337), Y => n791);
   U1239 : OAI211xp5_ASAP7_75t_R port map( A1 => n185, A2 => n73, B => n792, C 
                           => n793, Y => crossbar_out(16));
   U1240 : AOI222xp33_ASAP7_75t_R port map( A1 => n71, A2 => crossbar_in(272), 
                           B1 => n65, B2 => crossbar_in(400), C1 => n59, C2 => 
                           crossbar_in(336), Y => n793);
   U1241 : OAI211xp5_ASAP7_75t_R port map( A1 => n186, A2 => n73, B => n794, C 
                           => n795, Y => crossbar_out(15));
   U1242 : AOI222xp33_ASAP7_75t_R port map( A1 => n71, A2 => crossbar_in(271), 
                           B1 => n65, B2 => crossbar_in(399), C1 => n59, C2 => 
                           crossbar_in(335), Y => n795);
   U1243 : OAI211xp5_ASAP7_75t_R port map( A1 => n187, A2 => n73, B => n796, C 
                           => n797, Y => crossbar_out(14));
   U1244 : AOI222xp33_ASAP7_75t_R port map( A1 => n71, A2 => crossbar_in(270), 
                           B1 => n65, B2 => crossbar_in(398), C1 => n59, C2 => 
                           crossbar_in(334), Y => n797);
   U1245 : OAI211xp5_ASAP7_75t_R port map( A1 => n188, A2 => n73, B => n798, C 
                           => n799, Y => crossbar_out(13));
   U1246 : AOI222xp33_ASAP7_75t_R port map( A1 => n71, A2 => crossbar_in(269), 
                           B1 => n65, B2 => crossbar_in(397), C1 => n59, C2 => 
                           crossbar_in(333), Y => n799);
   U1247 : OAI211xp5_ASAP7_75t_R port map( A1 => n189, A2 => n73, B => n800, C 
                           => n801, Y => crossbar_out(12));
   U1248 : AOI222xp33_ASAP7_75t_R port map( A1 => n72, A2 => crossbar_in(268), 
                           B1 => n66, B2 => crossbar_in(396), C1 => n60, C2 => 
                           crossbar_in(332), Y => n801);
   U1249 : OAI211xp5_ASAP7_75t_R port map( A1 => n190, A2 => n73, B => n802, C 
                           => n803, Y => crossbar_out(11));
   U1250 : AOI222xp33_ASAP7_75t_R port map( A1 => n72, A2 => crossbar_in(267), 
                           B1 => n66, B2 => crossbar_in(395), C1 => n60, C2 => 
                           crossbar_in(331), Y => n803);
   U1251 : OAI211xp5_ASAP7_75t_R port map( A1 => n191, A2 => n73, B => n804, C 
                           => n805, Y => crossbar_out(10));
   U1252 : AOI222xp33_ASAP7_75t_R port map( A1 => n72, A2 => crossbar_in(266), 
                           B1 => n66, B2 => crossbar_in(394), C1 => n60, C2 => 
                           crossbar_in(330), Y => n805);
   U1253 : OAI211xp5_ASAP7_75t_R port map( A1 => n201, A2 => n73, B => n806, C 
                           => n807, Y => crossbar_out(0));
   U1254 : AOI222xp33_ASAP7_75t_R port map( A1 => n72, A2 => crossbar_in(256), 
                           B1 => n66, B2 => crossbar_in(384), C1 => n60, C2 => 
                           crossbar_in(320), Y => n807);
   U1255 : NAND3xp33_ASAP7_75t_R port map( A => n912, B => n911, C => n164, Y 
                           => n674);
   U128 : HB1xp67_ASAP7_75t_R port map( A => n537, Y => n131);
   U129 : HB1xp67_ASAP7_75t_R port map( A => n537, Y => n128);
   U130 : HB1xp67_ASAP7_75t_R port map( A => n537, Y => n129);
   U132 : HB1xp67_ASAP7_75t_R port map( A => n537, Y => n130);
   U133 : HB1xp67_ASAP7_75t_R port map( A => n537, Y => n126);
   U135 : HB1xp67_ASAP7_75t_R port map( A => n537, Y => n127);
   U136 : INVx1_ASAP7_75t_R port map( A => n171, Y => n165);
   U137 : HB1xp67_ASAP7_75t_R port map( A => n541, Y => n113);
   U139 : HB1xp67_ASAP7_75t_R port map( A => n541, Y => n112);
   U140 : HB1xp67_ASAP7_75t_R port map( A => n541, Y => n111);
   U141 : HB1xp67_ASAP7_75t_R port map( A => n541, Y => n110);
   U206 : HB1xp67_ASAP7_75t_R port map( A => n541, Y => n109);
   U207 : HB1xp67_ASAP7_75t_R port map( A => n541, Y => n108);
   U208 : HB1xp67_ASAP7_75t_R port map( A => n542, Y => n107);
   U210 : HB1xp67_ASAP7_75t_R port map( A => n538, Y => n125);
   U211 : HB1xp67_ASAP7_75t_R port map( A => n609, Y => n89);
   U212 : HB1xp67_ASAP7_75t_R port map( A => n610, Y => n83);
   U213 : HB1xp67_ASAP7_75t_R port map( A => n538, Y => n124);
   U214 : HB1xp67_ASAP7_75t_R port map( A => n538, Y => n123);
   U215 : HB1xp67_ASAP7_75t_R port map( A => n538, Y => n122);
   U216 : HB1xp67_ASAP7_75t_R port map( A => n407, Y => n152);
   U217 : HB1xp67_ASAP7_75t_R port map( A => n407, Y => n151);
   U218 : HB1xp67_ASAP7_75t_R port map( A => n407, Y => n149);
   U219 : HB1xp67_ASAP7_75t_R port map( A => n538, Y => n121);
   U220 : HB1xp67_ASAP7_75t_R port map( A => n538, Y => n120);
   U221 : HB1xp67_ASAP7_75t_R port map( A => n407, Y => n150);
   U222 : HB1xp67_ASAP7_75t_R port map( A => n542, Y => n106);
   U223 : HB1xp67_ASAP7_75t_R port map( A => n542, Y => n105);
   U224 : HB1xp67_ASAP7_75t_R port map( A => n542, Y => n104);
   U225 : HB1xp67_ASAP7_75t_R port map( A => n407, Y => n153);
   U226 : HB1xp67_ASAP7_75t_R port map( A => n542, Y => n103);
   U227 : HB1xp67_ASAP7_75t_R port map( A => n542, Y => n102);
   U228 : HB1xp67_ASAP7_75t_R port map( A => n406, Y => n157);
   U229 : HB1xp67_ASAP7_75t_R port map( A => n406, Y => n156);
   U230 : HB1xp67_ASAP7_75t_R port map( A => n406, Y => n155);
   U231 : HB1xp67_ASAP7_75t_R port map( A => n406, Y => n154);
   U232 : HB1xp67_ASAP7_75t_R port map( A => n406, Y => n158);
   U233 : HB1xp67_ASAP7_75t_R port map( A => n609, Y => n88);
   U234 : HB1xp67_ASAP7_75t_R port map( A => n609, Y => n87);
   U235 : HB1xp67_ASAP7_75t_R port map( A => n609, Y => n86);
   U236 : HB1xp67_ASAP7_75t_R port map( A => n609, Y => n85);
   U237 : HB1xp67_ASAP7_75t_R port map( A => n609, Y => n84);
   U238 : HB1xp67_ASAP7_75t_R port map( A => n610, Y => n82);
   U239 : HB1xp67_ASAP7_75t_R port map( A => n610, Y => n81);
   U240 : HB1xp67_ASAP7_75t_R port map( A => n610, Y => n80);
   U241 : HB1xp67_ASAP7_75t_R port map( A => n610, Y => n79);
   U242 : HB1xp67_ASAP7_75t_R port map( A => n610, Y => n78);
   U243 : HB1xp67_ASAP7_75t_R port map( A => n606, Y => n101);
   U244 : HB1xp67_ASAP7_75t_R port map( A => n403, Y => n159);
   U245 : HB1xp67_ASAP7_75t_R port map( A => n403, Y => n160);
   U246 : HB1xp67_ASAP7_75t_R port map( A => n403, Y => n161);
   U247 : HB1xp67_ASAP7_75t_R port map( A => n403, Y => n162);
   U248 : HB1xp67_ASAP7_75t_R port map( A => n403, Y => n163);
   U249 : HB1xp67_ASAP7_75t_R port map( A => n606, Y => n100);
   U250 : HB1xp67_ASAP7_75t_R port map( A => n606, Y => n99);
   U251 : HB1xp67_ASAP7_75t_R port map( A => n606, Y => n98);
   U252 : HB1xp67_ASAP7_75t_R port map( A => n606, Y => n96);
   U253 : HB1xp67_ASAP7_75t_R port map( A => n606, Y => n97);
   U254 : HB1xp67_ASAP7_75t_R port map( A => n408, Y => n147);
   U255 : HB1xp67_ASAP7_75t_R port map( A => n408, Y => n146);
   U256 : HB1xp67_ASAP7_75t_R port map( A => n408, Y => n145);
   U257 : HB1xp67_ASAP7_75t_R port map( A => n408, Y => n144);
   U258 : HB1xp67_ASAP7_75t_R port map( A => n408, Y => n148);
   U259 : HB1xp67_ASAP7_75t_R port map( A => n409, Y => n143);
   U260 : HB1xp67_ASAP7_75t_R port map( A => n409, Y => n142);
   U261 : HB1xp67_ASAP7_75t_R port map( A => n409, Y => n141);
   U262 : HB1xp67_ASAP7_75t_R port map( A => n409, Y => n140);
   U263 : HB1xp67_ASAP7_75t_R port map( A => n409, Y => n139);
   U264 : HB1xp67_ASAP7_75t_R port map( A => n409, Y => n138);
   U265 : HB1xp67_ASAP7_75t_R port map( A => crossbar_ctrl(18), Y => n171);
   U266 : HB1xp67_ASAP7_75t_R port map( A => n910, Y => n42);
   U267 : HB1xp67_ASAP7_75t_R port map( A => n910, Y => n37);
   U268 : HB1xp67_ASAP7_75t_R port map( A => n910, Y => n38);
   U269 : HB1xp67_ASAP7_75t_R port map( A => n910, Y => n39);
   U270 : HB1xp67_ASAP7_75t_R port map( A => n910, Y => n40);
   U271 : HB1xp67_ASAP7_75t_R port map( A => n910, Y => n41);
   U272 : HB1xp67_ASAP7_75t_R port map( A => crossbar_ctrl(18), Y => n170);
   U273 : HB1xp67_ASAP7_75t_R port map( A => crossbar_ctrl(18), Y => n169);
   U274 : HB1xp67_ASAP7_75t_R port map( A => crossbar_ctrl(18), Y => n168);
   U275 : HB1xp67_ASAP7_75t_R port map( A => crossbar_ctrl(18), Y => n167);
   U276 : HB1xp67_ASAP7_75t_R port map( A => crossbar_ctrl(18), Y => n166);
   U277 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(0), Y => n164);
   U278 : NOR2xp33_ASAP7_75t_R port map( A => n902, B => n901, Y => n541);
   U279 : NOR2xp33_ASAP7_75t_R port map( A => n901, B => crossbar_ctrl(9), Y =>
                           n542);
   U280 : NOR2xp33_ASAP7_75t_R port map( A => n906, B => n907, Y => n609);
   U281 : NOR2xp33_ASAP7_75t_R port map( A => n906, B => crossbar_ctrl(3), Y =>
                           n610);
   U282 : NOR2xp33_ASAP7_75t_R port map( A => n897, B => n899, Y => n407);
   U283 : HB1xp67_ASAP7_75t_R port map( A => n410, Y => n137);
   U284 : NOR2xp33_ASAP7_75t_R port map( A => n898, B => n899, Y => n406);
   U285 : HB1xp67_ASAP7_75t_R port map( A => n410, Y => n132);
   U286 : HB1xp67_ASAP7_75t_R port map( A => n904, Y => n18);
   U287 : HB1xp67_ASAP7_75t_R port map( A => n410, Y => n136);
   U288 : HB1xp67_ASAP7_75t_R port map( A => n410, Y => n135);
   U289 : HB1xp67_ASAP7_75t_R port map( A => n410, Y => n134);
   U290 : HB1xp67_ASAP7_75t_R port map( A => n410, Y => n133);
   U291 : HB1xp67_ASAP7_75t_R port map( A => n903, Y => n12);
   U292 : NOR2xp33_ASAP7_75t_R port map( A => n897, B => crossbar_ctrl(15), Y 
                           => n408);
   U293 : NOR2xp33_ASAP7_75t_R port map( A => n898, B => crossbar_ctrl(15), Y 
                           => n409);
   U294 : HB1xp67_ASAP7_75t_R port map( A => n903, Y => n7);
   U295 : HB1xp67_ASAP7_75t_R port map( A => n903, Y => n8);
   U296 : HB1xp67_ASAP7_75t_R port map( A => n903, Y => n9);
   U297 : HB1xp67_ASAP7_75t_R port map( A => n903, Y => n10);
   U298 : HB1xp67_ASAP7_75t_R port map( A => n903, Y => n11);
   U299 : HB1xp67_ASAP7_75t_R port map( A => n904, Y => n13);
   U300 : HB1xp67_ASAP7_75t_R port map( A => n904, Y => n14);
   U301 : HB1xp67_ASAP7_75t_R port map( A => n904, Y => n15);
   U302 : HB1xp67_ASAP7_75t_R port map( A => n904, Y => n16);
   U303 : HB1xp67_ASAP7_75t_R port map( A => n904, Y => n17);
   U304 : HB1xp67_ASAP7_75t_R port map( A => n540, Y => n119);
   U305 : HB1xp67_ASAP7_75t_R port map( A => n540, Y => n118);
   U306 : HB1xp67_ASAP7_75t_R port map( A => n540, Y => n117);
   U307 : HB1xp67_ASAP7_75t_R port map( A => n540, Y => n116);
   U308 : HB1xp67_ASAP7_75t_R port map( A => n540, Y => n115);
   U309 : HB1xp67_ASAP7_75t_R port map( A => n540, Y => n114);
   U310 : HB1xp67_ASAP7_75t_R port map( A => n608, Y => n95);
   U311 : NOR3xp33_ASAP7_75t_R port map( A => crossbar_ctrl(16), B => 
                           crossbar_ctrl(17), C => n899, Y => n410);
   U312 : HB1xp67_ASAP7_75t_R port map( A => n608, Y => n90);
   U313 : HB1xp67_ASAP7_75t_R port map( A => n608, Y => n94);
   U314 : HB1xp67_ASAP7_75t_R port map( A => n608, Y => n93);
   U315 : HB1xp67_ASAP7_75t_R port map( A => n608, Y => n92);
   U316 : HB1xp67_ASAP7_75t_R port map( A => n608, Y => n91);
   U317 : HB1xp67_ASAP7_75t_R port map( A => n900, Y => n6);
   U318 : HB1xp67_ASAP7_75t_R port map( A => n900, Y => n1);
   U319 : HB1xp67_ASAP7_75t_R port map( A => n900, Y => n2);
   U320 : HB1xp67_ASAP7_75t_R port map( A => n900, Y => n3);
   U321 : HB1xp67_ASAP7_75t_R port map( A => n900, Y => n4);
   U322 : HB1xp67_ASAP7_75t_R port map( A => n900, Y => n5);
   U323 : HB1xp67_ASAP7_75t_R port map( A => n905, Y => n24);
   U324 : HB1xp67_ASAP7_75t_R port map( A => n905, Y => n19);
   U325 : HB1xp67_ASAP7_75t_R port map( A => n905, Y => n20);
   U326 : HB1xp67_ASAP7_75t_R port map( A => n905, Y => n21);
   U327 : HB1xp67_ASAP7_75t_R port map( A => n905, Y => n23);
   U328 : HB1xp67_ASAP7_75t_R port map( A => n905, Y => n22);
   U329 : HB1xp67_ASAP7_75t_R port map( A => n909, Y => n36);
   U330 : HB1xp67_ASAP7_75t_R port map( A => n908, Y => n30);
   U331 : HB1xp67_ASAP7_75t_R port map( A => n909, Y => n31);
   U332 : HB1xp67_ASAP7_75t_R port map( A => n909, Y => n32);
   U333 : HB1xp67_ASAP7_75t_R port map( A => n909, Y => n33);
   U334 : HB1xp67_ASAP7_75t_R port map( A => n909, Y => n34);
   U335 : HB1xp67_ASAP7_75t_R port map( A => n909, Y => n35);
   U336 : HB1xp67_ASAP7_75t_R port map( A => n908, Y => n25);
   U337 : HB1xp67_ASAP7_75t_R port map( A => n908, Y => n26);
   U338 : HB1xp67_ASAP7_75t_R port map( A => n908, Y => n27);
   U339 : HB1xp67_ASAP7_75t_R port map( A => n908, Y => n28);
   U340 : HB1xp67_ASAP7_75t_R port map( A => n908, Y => n29);
   U341 : HB1xp67_ASAP7_75t_R port map( A => n678, Y => n66);
   U342 : HB1xp67_ASAP7_75t_R port map( A => n677, Y => n72);
   U343 : HB1xp67_ASAP7_75t_R port map( A => n674, Y => n73);
   U344 : HB1xp67_ASAP7_75t_R port map( A => n674, Y => n74);
   U345 : HB1xp67_ASAP7_75t_R port map( A => n674, Y => n75);
   U346 : HB1xp67_ASAP7_75t_R port map( A => n674, Y => n76);
   U347 : HB1xp67_ASAP7_75t_R port map( A => n679, Y => n60);
   U348 : HB1xp67_ASAP7_75t_R port map( A => n674, Y => n77);
   U349 : HB1xp67_ASAP7_75t_R port map( A => n678, Y => n65);
   U350 : HB1xp67_ASAP7_75t_R port map( A => n678, Y => n64);
   U351 : HB1xp67_ASAP7_75t_R port map( A => n678, Y => n63);
   U352 : HB1xp67_ASAP7_75t_R port map( A => n678, Y => n62);
   U353 : HB1xp67_ASAP7_75t_R port map( A => n678, Y => n61);
   U354 : HB1xp67_ASAP7_75t_R port map( A => n677, Y => n71);
   U355 : HB1xp67_ASAP7_75t_R port map( A => n677, Y => n70);
   U356 : HB1xp67_ASAP7_75t_R port map( A => n677, Y => n69);
   U357 : HB1xp67_ASAP7_75t_R port map( A => n677, Y => n68);
   U358 : HB1xp67_ASAP7_75t_R port map( A => n677, Y => n67);
   U359 : HB1xp67_ASAP7_75t_R port map( A => n679, Y => n59);
   U360 : HB1xp67_ASAP7_75t_R port map( A => n679, Y => n58);
   U361 : HB1xp67_ASAP7_75t_R port map( A => n679, Y => n57);
   U362 : HB1xp67_ASAP7_75t_R port map( A => n679, Y => n56);
   U363 : HB1xp67_ASAP7_75t_R port map( A => n679, Y => n55);
   U364 : HB1xp67_ASAP7_75t_R port map( A => n680, Y => n54);
   U365 : HB1xp67_ASAP7_75t_R port map( A => n680, Y => n53);
   U366 : HB1xp67_ASAP7_75t_R port map( A => n680, Y => n52);
   U367 : HB1xp67_ASAP7_75t_R port map( A => n680, Y => n51);
   U368 : HB1xp67_ASAP7_75t_R port map( A => n680, Y => n50);
   U369 : HB1xp67_ASAP7_75t_R port map( A => n680, Y => n49);
   U370 : NOR3xp33_ASAP7_75t_R port map( A => crossbar_ctrl(10), B => 
                           crossbar_ctrl(11), C => n902, Y => n540);
   U371 : NOR3xp33_ASAP7_75t_R port map( A => crossbar_ctrl(4), B => 
                           crossbar_ctrl(5), C => n907, Y => n608);
   U372 : NOR2xp33_ASAP7_75t_R port map( A => n911, B => n164, Y => n678);
   U373 : HB1xp67_ASAP7_75t_R port map( A => n681, Y => n48);
   U374 : NOR2xp33_ASAP7_75t_R port map( A => n912, B => n164, Y => n677);
   U375 : NOR2xp33_ASAP7_75t_R port map( A => n911, B => crossbar_ctrl(0), Y =>
                           n679);
   U376 : HB1xp67_ASAP7_75t_R port map( A => n681, Y => n47);
   U377 : HB1xp67_ASAP7_75t_R port map( A => n681, Y => n46);
   U378 : HB1xp67_ASAP7_75t_R port map( A => n681, Y => n45);
   U379 : HB1xp67_ASAP7_75t_R port map( A => n681, Y => n44);
   U380 : HB1xp67_ASAP7_75t_R port map( A => n681, Y => n43);
   U381 : NOR2xp33_ASAP7_75t_R port map( A => n912, B => crossbar_ctrl(0), Y =>
                           n680);
   U382 : NOR3xp33_ASAP7_75t_R port map( A => crossbar_ctrl(1), B => 
                           crossbar_ctrl(2), C => n164, Y => n681);
   U383 : INVx1_ASAP7_75t_R port map( A => crossbar_in(93), Y => n172);
   U384 : INVx1_ASAP7_75t_R port map( A => crossbar_in(92), Y => n173);
   U385 : INVx1_ASAP7_75t_R port map( A => crossbar_in(91), Y => n174);
   U386 : INVx1_ASAP7_75t_R port map( A => crossbar_in(90), Y => n175);
   U387 : INVx1_ASAP7_75t_R port map( A => crossbar_in(89), Y => n176);
   U388 : INVx1_ASAP7_75t_R port map( A => crossbar_in(88), Y => n177);
   U389 : INVx1_ASAP7_75t_R port map( A => crossbar_in(87), Y => n178);
   U390 : INVx1_ASAP7_75t_R port map( A => crossbar_in(86), Y => n179);
   U391 : INVx1_ASAP7_75t_R port map( A => crossbar_in(85), Y => n180);
   U392 : INVx1_ASAP7_75t_R port map( A => crossbar_in(84), Y => n181);
   U393 : INVx1_ASAP7_75t_R port map( A => crossbar_in(83), Y => n182);
   U394 : INVx1_ASAP7_75t_R port map( A => crossbar_in(82), Y => n183);
   U395 : INVx1_ASAP7_75t_R port map( A => crossbar_in(81), Y => n184);
   U396 : INVx1_ASAP7_75t_R port map( A => crossbar_in(80), Y => n185);
   U397 : INVx1_ASAP7_75t_R port map( A => crossbar_in(79), Y => n186);
   U398 : INVx1_ASAP7_75t_R port map( A => crossbar_in(78), Y => n187);
   U399 : INVx1_ASAP7_75t_R port map( A => crossbar_in(77), Y => n188);
   U400 : INVx1_ASAP7_75t_R port map( A => crossbar_in(76), Y => n189);
   U401 : INVx1_ASAP7_75t_R port map( A => crossbar_in(75), Y => n190);
   U402 : INVx1_ASAP7_75t_R port map( A => crossbar_in(74), Y => n191);
   U403 : INVx1_ASAP7_75t_R port map( A => crossbar_in(73), Y => n192);
   U404 : INVx1_ASAP7_75t_R port map( A => crossbar_in(72), Y => n193);
   U405 : INVx1_ASAP7_75t_R port map( A => crossbar_in(71), Y => n194);
   U406 : INVx1_ASAP7_75t_R port map( A => crossbar_in(70), Y => n195);
   U407 : INVx1_ASAP7_75t_R port map( A => crossbar_in(69), Y => n196);
   U408 : INVx1_ASAP7_75t_R port map( A => crossbar_in(68), Y => n197);
   U409 : INVx1_ASAP7_75t_R port map( A => crossbar_in(67), Y => n198);
   U410 : INVx1_ASAP7_75t_R port map( A => crossbar_in(66), Y => n199);
   U411 : INVx1_ASAP7_75t_R port map( A => crossbar_in(65), Y => n200);
   U412 : INVx1_ASAP7_75t_R port map( A => crossbar_in(64), Y => n201);
   U413 : INVx1_ASAP7_75t_R port map( A => crossbar_in(127), Y => n202);
   U414 : INVx1_ASAP7_75t_R port map( A => crossbar_in(126), Y => n203);
   U415 : INVx1_ASAP7_75t_R port map( A => crossbar_in(125), Y => n204);
   U416 : INVx1_ASAP7_75t_R port map( A => crossbar_in(124), Y => n205);
   U417 : INVx1_ASAP7_75t_R port map( A => crossbar_in(123), Y => n206);
   U418 : INVx1_ASAP7_75t_R port map( A => crossbar_in(122), Y => n207);
   U419 : INVx1_ASAP7_75t_R port map( A => crossbar_in(121), Y => n208);
   U420 : INVx1_ASAP7_75t_R port map( A => crossbar_in(120), Y => n209);
   U421 : INVx1_ASAP7_75t_R port map( A => crossbar_in(119), Y => n210);
   U422 : INVx1_ASAP7_75t_R port map( A => crossbar_in(118), Y => n211);
   U423 : INVx1_ASAP7_75t_R port map( A => crossbar_in(117), Y => n212);
   U424 : INVx1_ASAP7_75t_R port map( A => crossbar_in(116), Y => n213);
   U425 : INVx1_ASAP7_75t_R port map( A => crossbar_in(115), Y => n214);
   U426 : INVx1_ASAP7_75t_R port map( A => crossbar_in(114), Y => n215);
   U427 : INVx1_ASAP7_75t_R port map( A => crossbar_in(113), Y => n216);
   U428 : INVx1_ASAP7_75t_R port map( A => crossbar_in(112), Y => n217);
   U429 : INVx1_ASAP7_75t_R port map( A => crossbar_in(111), Y => n218);
   U430 : INVx1_ASAP7_75t_R port map( A => crossbar_in(110), Y => n219);
   U431 : INVx1_ASAP7_75t_R port map( A => crossbar_in(109), Y => n220);
   U432 : INVx1_ASAP7_75t_R port map( A => crossbar_in(108), Y => n221);
   U433 : INVx1_ASAP7_75t_R port map( A => crossbar_in(107), Y => n222);
   U434 : INVx1_ASAP7_75t_R port map( A => crossbar_in(106), Y => n223);
   U435 : INVx1_ASAP7_75t_R port map( A => crossbar_in(105), Y => n224);
   U436 : INVx1_ASAP7_75t_R port map( A => crossbar_in(104), Y => n225);
   U437 : INVx1_ASAP7_75t_R port map( A => crossbar_in(103), Y => n226);
   U438 : INVx1_ASAP7_75t_R port map( A => crossbar_in(102), Y => n227);
   U439 : INVx1_ASAP7_75t_R port map( A => crossbar_in(101), Y => n228);
   U440 : INVx1_ASAP7_75t_R port map( A => crossbar_in(100), Y => n229);
   U441 : INVx1_ASAP7_75t_R port map( A => crossbar_in(99), Y => n230);
   U442 : INVx1_ASAP7_75t_R port map( A => crossbar_in(98), Y => n231);
   U443 : INVx1_ASAP7_75t_R port map( A => crossbar_in(97), Y => n232);
   U444 : INVx1_ASAP7_75t_R port map( A => crossbar_in(96), Y => n233);
   U445 : INVx1_ASAP7_75t_R port map( A => crossbar_in(95), Y => n234);
   U446 : INVx1_ASAP7_75t_R port map( A => crossbar_in(94), Y => n235);
   U447 : INVx1_ASAP7_75t_R port map( A => crossbar_in(285), Y => n236);
   U448 : INVx1_ASAP7_75t_R port map( A => crossbar_in(284), Y => n237);
   U449 : INVx1_ASAP7_75t_R port map( A => crossbar_in(283), Y => n238);
   U450 : INVx1_ASAP7_75t_R port map( A => crossbar_in(282), Y => n239);
   U451 : INVx1_ASAP7_75t_R port map( A => crossbar_in(281), Y => n240);
   U452 : INVx1_ASAP7_75t_R port map( A => crossbar_in(280), Y => n241);
   U453 : INVx1_ASAP7_75t_R port map( A => crossbar_in(279), Y => n242);
   U454 : INVx1_ASAP7_75t_R port map( A => crossbar_in(278), Y => n243);
   U455 : INVx1_ASAP7_75t_R port map( A => crossbar_in(277), Y => n244);
   U456 : INVx1_ASAP7_75t_R port map( A => crossbar_in(276), Y => n245);
   U457 : INVx1_ASAP7_75t_R port map( A => crossbar_in(275), Y => n246);
   U458 : INVx1_ASAP7_75t_R port map( A => crossbar_in(274), Y => n247);
   U459 : INVx1_ASAP7_75t_R port map( A => crossbar_in(273), Y => n248);
   U460 : INVx1_ASAP7_75t_R port map( A => crossbar_in(272), Y => n249);
   U461 : INVx1_ASAP7_75t_R port map( A => crossbar_in(271), Y => n250);
   U462 : INVx1_ASAP7_75t_R port map( A => crossbar_in(270), Y => n251);
   U463 : INVx1_ASAP7_75t_R port map( A => crossbar_in(269), Y => n252);
   U464 : INVx1_ASAP7_75t_R port map( A => crossbar_in(268), Y => n253);
   U465 : INVx1_ASAP7_75t_R port map( A => crossbar_in(267), Y => n254);
   U466 : INVx1_ASAP7_75t_R port map( A => crossbar_in(266), Y => n255);
   U467 : INVx1_ASAP7_75t_R port map( A => crossbar_in(265), Y => n256);
   U468 : INVx1_ASAP7_75t_R port map( A => crossbar_in(264), Y => n257);
   U469 : INVx1_ASAP7_75t_R port map( A => crossbar_in(263), Y => n258);
   U470 : INVx1_ASAP7_75t_R port map( A => crossbar_in(262), Y => n259);
   U471 : INVx1_ASAP7_75t_R port map( A => crossbar_in(261), Y => n260);
   U472 : INVx1_ASAP7_75t_R port map( A => crossbar_in(260), Y => n261);
   U473 : INVx1_ASAP7_75t_R port map( A => crossbar_in(259), Y => n262);
   U474 : INVx1_ASAP7_75t_R port map( A => crossbar_in(258), Y => n263);
   U475 : INVx1_ASAP7_75t_R port map( A => crossbar_in(257), Y => n264);
   U476 : INVx1_ASAP7_75t_R port map( A => crossbar_in(256), Y => n265);
   U477 : INVx1_ASAP7_75t_R port map( A => crossbar_in(319), Y => n266);
   U478 : INVx1_ASAP7_75t_R port map( A => crossbar_in(318), Y => n267);
   U479 : INVx1_ASAP7_75t_R port map( A => crossbar_in(317), Y => n268);
   U480 : INVx1_ASAP7_75t_R port map( A => crossbar_in(316), Y => n269);
   U481 : INVx1_ASAP7_75t_R port map( A => crossbar_in(315), Y => n270);
   U482 : INVx1_ASAP7_75t_R port map( A => crossbar_in(314), Y => n271);
   U483 : INVx1_ASAP7_75t_R port map( A => crossbar_in(313), Y => n272);
   U484 : INVx1_ASAP7_75t_R port map( A => crossbar_in(312), Y => n273);
   U485 : INVx1_ASAP7_75t_R port map( A => crossbar_in(311), Y => n274);
   U486 : INVx1_ASAP7_75t_R port map( A => crossbar_in(310), Y => n275);
   U487 : INVx1_ASAP7_75t_R port map( A => crossbar_in(309), Y => n276);
   U488 : INVx1_ASAP7_75t_R port map( A => crossbar_in(308), Y => n277);
   U489 : INVx1_ASAP7_75t_R port map( A => crossbar_in(307), Y => n278);
   U490 : INVx1_ASAP7_75t_R port map( A => crossbar_in(306), Y => n279);
   U491 : INVx1_ASAP7_75t_R port map( A => crossbar_in(305), Y => n280);
   U492 : INVx1_ASAP7_75t_R port map( A => crossbar_in(304), Y => n281);
   U493 : INVx1_ASAP7_75t_R port map( A => crossbar_in(303), Y => n282);
   U494 : INVx1_ASAP7_75t_R port map( A => crossbar_in(302), Y => n283);
   U495 : INVx1_ASAP7_75t_R port map( A => crossbar_in(301), Y => n284);
   U496 : INVx1_ASAP7_75t_R port map( A => crossbar_in(300), Y => n285);
   U497 : INVx1_ASAP7_75t_R port map( A => crossbar_in(299), Y => n286);
   U498 : INVx1_ASAP7_75t_R port map( A => crossbar_in(298), Y => n287);
   U499 : INVx1_ASAP7_75t_R port map( A => crossbar_in(297), Y => n288);
   U500 : INVx1_ASAP7_75t_R port map( A => crossbar_in(296), Y => n289);
   U501 : INVx1_ASAP7_75t_R port map( A => crossbar_in(295), Y => n290);
   U502 : INVx1_ASAP7_75t_R port map( A => crossbar_in(294), Y => n291);
   U503 : INVx1_ASAP7_75t_R port map( A => crossbar_in(293), Y => n292);
   U504 : INVx1_ASAP7_75t_R port map( A => crossbar_in(292), Y => n293);
   U505 : INVx1_ASAP7_75t_R port map( A => crossbar_in(291), Y => n294);
   U506 : INVx1_ASAP7_75t_R port map( A => crossbar_in(290), Y => n295);
   U507 : INVx1_ASAP7_75t_R port map( A => crossbar_in(289), Y => n296);
   U508 : INVx1_ASAP7_75t_R port map( A => crossbar_in(288), Y => n297);
   U509 : INVx1_ASAP7_75t_R port map( A => crossbar_in(287), Y => n298);
   U510 : INVx1_ASAP7_75t_R port map( A => crossbar_in(286), Y => n299);
   U511 : INVx1_ASAP7_75t_R port map( A => crossbar_in(349), Y => n300);
   U512 : INVx1_ASAP7_75t_R port map( A => crossbar_in(348), Y => n301);
   U513 : INVx1_ASAP7_75t_R port map( A => crossbar_in(347), Y => n302);
   U514 : INVx1_ASAP7_75t_R port map( A => crossbar_in(346), Y => n303);
   U515 : INVx1_ASAP7_75t_R port map( A => crossbar_in(345), Y => n304);
   U516 : INVx1_ASAP7_75t_R port map( A => crossbar_in(344), Y => n305);
   U517 : INVx1_ASAP7_75t_R port map( A => crossbar_in(343), Y => n306);
   U518 : INVx1_ASAP7_75t_R port map( A => crossbar_in(342), Y => n307);
   U519 : INVx1_ASAP7_75t_R port map( A => crossbar_in(341), Y => n308);
   U520 : INVx1_ASAP7_75t_R port map( A => crossbar_in(340), Y => n309);
   U521 : INVx1_ASAP7_75t_R port map( A => crossbar_in(339), Y => n310);
   U522 : INVx1_ASAP7_75t_R port map( A => crossbar_in(338), Y => n311);
   U523 : INVx1_ASAP7_75t_R port map( A => crossbar_in(337), Y => n312);
   U524 : INVx1_ASAP7_75t_R port map( A => crossbar_in(336), Y => n313);
   U525 : INVx1_ASAP7_75t_R port map( A => crossbar_in(335), Y => n314);
   U526 : INVx1_ASAP7_75t_R port map( A => crossbar_in(334), Y => n315);
   U527 : INVx1_ASAP7_75t_R port map( A => crossbar_in(333), Y => n316);
   U528 : INVx1_ASAP7_75t_R port map( A => crossbar_in(332), Y => n317);
   U529 : INVx1_ASAP7_75t_R port map( A => crossbar_in(331), Y => n318);
   U530 : INVx1_ASAP7_75t_R port map( A => crossbar_in(330), Y => n319);
   U531 : INVx1_ASAP7_75t_R port map( A => crossbar_in(329), Y => n320);
   U532 : INVx1_ASAP7_75t_R port map( A => crossbar_in(328), Y => n321);
   U533 : INVx1_ASAP7_75t_R port map( A => crossbar_in(327), Y => n322);
   U534 : INVx1_ASAP7_75t_R port map( A => crossbar_in(326), Y => n323);
   U535 : INVx1_ASAP7_75t_R port map( A => crossbar_in(325), Y => n324);
   U536 : INVx1_ASAP7_75t_R port map( A => crossbar_in(324), Y => n325);
   U537 : INVx1_ASAP7_75t_R port map( A => crossbar_in(323), Y => n326);
   U538 : INVx1_ASAP7_75t_R port map( A => crossbar_in(322), Y => n327);
   U539 : INVx1_ASAP7_75t_R port map( A => crossbar_in(321), Y => n328);
   U540 : INVx1_ASAP7_75t_R port map( A => crossbar_in(320), Y => n329);
   U541 : INVx1_ASAP7_75t_R port map( A => crossbar_in(383), Y => n330);
   U542 : INVx1_ASAP7_75t_R port map( A => crossbar_in(382), Y => n331);
   U543 : INVx1_ASAP7_75t_R port map( A => crossbar_in(381), Y => n332);
   U544 : INVx1_ASAP7_75t_R port map( A => crossbar_in(380), Y => n333);
   U545 : INVx1_ASAP7_75t_R port map( A => crossbar_in(379), Y => n334);
   U546 : INVx1_ASAP7_75t_R port map( A => crossbar_in(378), Y => n335);
   U547 : INVx1_ASAP7_75t_R port map( A => crossbar_in(377), Y => n336);
   U548 : INVx1_ASAP7_75t_R port map( A => crossbar_in(376), Y => n337);
   U549 : INVx1_ASAP7_75t_R port map( A => crossbar_in(375), Y => n338);
   U550 : INVx1_ASAP7_75t_R port map( A => crossbar_in(374), Y => n339);
   U551 : INVx1_ASAP7_75t_R port map( A => crossbar_in(373), Y => n340);
   U552 : INVx1_ASAP7_75t_R port map( A => crossbar_in(372), Y => n341);
   U553 : INVx1_ASAP7_75t_R port map( A => crossbar_in(371), Y => n342);
   U554 : INVx1_ASAP7_75t_R port map( A => crossbar_in(370), Y => n343);
   U555 : INVx1_ASAP7_75t_R port map( A => crossbar_in(369), Y => n344);
   U556 : INVx1_ASAP7_75t_R port map( A => crossbar_in(368), Y => n345);
   U557 : INVx1_ASAP7_75t_R port map( A => crossbar_in(367), Y => n346);
   U558 : INVx1_ASAP7_75t_R port map( A => crossbar_in(366), Y => n347);
   U559 : INVx1_ASAP7_75t_R port map( A => crossbar_in(365), Y => n348);
   U560 : INVx1_ASAP7_75t_R port map( A => crossbar_in(364), Y => n349);
   U561 : INVx1_ASAP7_75t_R port map( A => crossbar_in(363), Y => n350);
   U562 : INVx1_ASAP7_75t_R port map( A => crossbar_in(362), Y => n351);
   U563 : INVx1_ASAP7_75t_R port map( A => crossbar_in(361), Y => n352);
   U564 : INVx1_ASAP7_75t_R port map( A => crossbar_in(360), Y => n353);
   U565 : INVx1_ASAP7_75t_R port map( A => crossbar_in(359), Y => n354);
   U566 : INVx1_ASAP7_75t_R port map( A => crossbar_in(358), Y => n355);
   U567 : INVx1_ASAP7_75t_R port map( A => crossbar_in(357), Y => n356);
   U568 : INVx1_ASAP7_75t_R port map( A => crossbar_in(356), Y => n357);
   U569 : INVx1_ASAP7_75t_R port map( A => crossbar_in(355), Y => n358);
   U570 : INVx1_ASAP7_75t_R port map( A => crossbar_in(354), Y => n359);
   U571 : INVx1_ASAP7_75t_R port map( A => crossbar_in(353), Y => n360);
   U572 : INVx1_ASAP7_75t_R port map( A => crossbar_in(352), Y => n361);
   U573 : INVx1_ASAP7_75t_R port map( A => crossbar_in(351), Y => n362);
   U574 : INVx1_ASAP7_75t_R port map( A => crossbar_in(350), Y => n363);
   U575 : INVx1_ASAP7_75t_R port map( A => crossbar_in(413), Y => n364);
   U576 : INVx1_ASAP7_75t_R port map( A => crossbar_in(412), Y => n365);
   U577 : INVx1_ASAP7_75t_R port map( A => crossbar_in(411), Y => n366);
   U578 : INVx1_ASAP7_75t_R port map( A => crossbar_in(410), Y => n367);
   U579 : INVx1_ASAP7_75t_R port map( A => crossbar_in(409), Y => n368);
   U580 : INVx1_ASAP7_75t_R port map( A => crossbar_in(408), Y => n369);
   U581 : INVx1_ASAP7_75t_R port map( A => crossbar_in(407), Y => n370);
   U582 : INVx1_ASAP7_75t_R port map( A => crossbar_in(406), Y => n371);
   U583 : INVx1_ASAP7_75t_R port map( A => crossbar_in(405), Y => n372);
   U584 : INVx1_ASAP7_75t_R port map( A => crossbar_in(404), Y => n373);
   U585 : INVx1_ASAP7_75t_R port map( A => crossbar_in(403), Y => n374);
   U586 : INVx1_ASAP7_75t_R port map( A => crossbar_in(402), Y => n375);
   U587 : INVx1_ASAP7_75t_R port map( A => crossbar_in(401), Y => n376);
   U588 : INVx1_ASAP7_75t_R port map( A => crossbar_in(400), Y => n377);
   U589 : INVx1_ASAP7_75t_R port map( A => crossbar_in(399), Y => n378);
   U590 : INVx1_ASAP7_75t_R port map( A => crossbar_in(398), Y => n379);
   U591 : INVx1_ASAP7_75t_R port map( A => crossbar_in(397), Y => n380);
   U592 : INVx1_ASAP7_75t_R port map( A => crossbar_in(396), Y => n381);
   U593 : INVx1_ASAP7_75t_R port map( A => crossbar_in(395), Y => n382);
   U594 : INVx1_ASAP7_75t_R port map( A => crossbar_in(394), Y => n383);
   U595 : INVx1_ASAP7_75t_R port map( A => crossbar_in(393), Y => n384);
   U596 : INVx1_ASAP7_75t_R port map( A => crossbar_in(392), Y => n385);
   U597 : INVx1_ASAP7_75t_R port map( A => crossbar_in(391), Y => n386);
   U598 : INVx1_ASAP7_75t_R port map( A => crossbar_in(390), Y => n387);
   U599 : INVx1_ASAP7_75t_R port map( A => crossbar_in(389), Y => n388);
   U600 : INVx1_ASAP7_75t_R port map( A => crossbar_in(388), Y => n389);
   U601 : INVx1_ASAP7_75t_R port map( A => crossbar_in(387), Y => n390);
   U602 : INVx1_ASAP7_75t_R port map( A => crossbar_in(386), Y => n391);
   U603 : INVx1_ASAP7_75t_R port map( A => crossbar_in(385), Y => n392);
   U604 : INVx1_ASAP7_75t_R port map( A => crossbar_in(384), Y => n393);
   U605 : INVx1_ASAP7_75t_R port map( A => crossbar_in(447), Y => n394);
   U606 : INVx1_ASAP7_75t_R port map( A => crossbar_in(446), Y => n395);
   U607 : INVx1_ASAP7_75t_R port map( A => crossbar_in(445), Y => n396);
   U608 : INVx1_ASAP7_75t_R port map( A => crossbar_in(444), Y => n397);
   U609 : INVx1_ASAP7_75t_R port map( A => crossbar_in(443), Y => n398);
   U610 : INVx1_ASAP7_75t_R port map( A => crossbar_in(442), Y => n399);
   U611 : INVx1_ASAP7_75t_R port map( A => crossbar_in(441), Y => n400);
   U612 : INVx1_ASAP7_75t_R port map( A => crossbar_in(440), Y => n401);
   U613 : INVx1_ASAP7_75t_R port map( A => crossbar_in(439), Y => n402);
   U1256 : INVx1_ASAP7_75t_R port map( A => crossbar_in(438), Y => n808);
   U1257 : INVx1_ASAP7_75t_R port map( A => crossbar_in(437), Y => n809);
   U1258 : INVx1_ASAP7_75t_R port map( A => crossbar_in(436), Y => n810);
   U1259 : INVx1_ASAP7_75t_R port map( A => crossbar_in(435), Y => n811);
   U1260 : INVx1_ASAP7_75t_R port map( A => crossbar_in(434), Y => n812);
   U1261 : INVx1_ASAP7_75t_R port map( A => crossbar_in(433), Y => n813);
   U1262 : INVx1_ASAP7_75t_R port map( A => crossbar_in(432), Y => n814);
   U1263 : INVx1_ASAP7_75t_R port map( A => crossbar_in(431), Y => n815);
   U1264 : INVx1_ASAP7_75t_R port map( A => crossbar_in(430), Y => n816);
   U1265 : INVx1_ASAP7_75t_R port map( A => crossbar_in(429), Y => n817);
   U1266 : INVx1_ASAP7_75t_R port map( A => crossbar_in(428), Y => n818);
   U1267 : INVx1_ASAP7_75t_R port map( A => crossbar_in(427), Y => n819);
   U1268 : INVx1_ASAP7_75t_R port map( A => crossbar_in(426), Y => n820);
   U1269 : INVx1_ASAP7_75t_R port map( A => crossbar_in(425), Y => n821);
   U1270 : INVx1_ASAP7_75t_R port map( A => crossbar_in(424), Y => n822);
   U1271 : INVx1_ASAP7_75t_R port map( A => crossbar_in(423), Y => n823);
   U1272 : INVx1_ASAP7_75t_R port map( A => crossbar_in(422), Y => n824);
   U1273 : INVx1_ASAP7_75t_R port map( A => crossbar_in(421), Y => n825);
   U1274 : INVx1_ASAP7_75t_R port map( A => crossbar_in(420), Y => n826);
   U1275 : INVx1_ASAP7_75t_R port map( A => crossbar_in(419), Y => n827);
   U1276 : INVx1_ASAP7_75t_R port map( A => crossbar_in(418), Y => n828);
   U1277 : INVx1_ASAP7_75t_R port map( A => crossbar_in(417), Y => n829);
   U1278 : INVx1_ASAP7_75t_R port map( A => crossbar_in(416), Y => n830);
   U1279 : INVx1_ASAP7_75t_R port map( A => crossbar_in(415), Y => n831);
   U1280 : INVx1_ASAP7_75t_R port map( A => crossbar_in(414), Y => n832);
   U1281 : INVx1_ASAP7_75t_R port map( A => crossbar_in(157), Y => n833);
   U1282 : INVx1_ASAP7_75t_R port map( A => crossbar_in(156), Y => n834);
   U1283 : INVx1_ASAP7_75t_R port map( A => crossbar_in(155), Y => n835);
   U1284 : INVx1_ASAP7_75t_R port map( A => crossbar_in(154), Y => n836);
   U1285 : INVx1_ASAP7_75t_R port map( A => crossbar_in(153), Y => n837);
   U1286 : INVx1_ASAP7_75t_R port map( A => crossbar_in(152), Y => n838);
   U1287 : INVx1_ASAP7_75t_R port map( A => crossbar_in(151), Y => n839);
   U1288 : INVx1_ASAP7_75t_R port map( A => crossbar_in(150), Y => n840);
   U1289 : INVx1_ASAP7_75t_R port map( A => crossbar_in(149), Y => n841);
   U1290 : INVx1_ASAP7_75t_R port map( A => crossbar_in(148), Y => n842);
   U1291 : INVx1_ASAP7_75t_R port map( A => crossbar_in(147), Y => n843);
   U1292 : INVx1_ASAP7_75t_R port map( A => crossbar_in(146), Y => n844);
   U1293 : INVx1_ASAP7_75t_R port map( A => crossbar_in(145), Y => n845);
   U1294 : INVx1_ASAP7_75t_R port map( A => crossbar_in(144), Y => n846);
   U1295 : INVx1_ASAP7_75t_R port map( A => crossbar_in(143), Y => n847);
   U1296 : INVx1_ASAP7_75t_R port map( A => crossbar_in(142), Y => n848);
   U1297 : INVx1_ASAP7_75t_R port map( A => crossbar_in(141), Y => n849);
   U1298 : INVx1_ASAP7_75t_R port map( A => crossbar_in(140), Y => n850);
   U1299 : INVx1_ASAP7_75t_R port map( A => crossbar_in(139), Y => n851);
   U1300 : INVx1_ASAP7_75t_R port map( A => crossbar_in(138), Y => n852);
   U1301 : INVx1_ASAP7_75t_R port map( A => crossbar_in(137), Y => n853);
   U1302 : INVx1_ASAP7_75t_R port map( A => crossbar_in(136), Y => n854);
   U1303 : INVx1_ASAP7_75t_R port map( A => crossbar_in(135), Y => n855);
   U1304 : INVx1_ASAP7_75t_R port map( A => crossbar_in(134), Y => n856);
   U1305 : INVx1_ASAP7_75t_R port map( A => crossbar_in(133), Y => n857);
   U1306 : INVx1_ASAP7_75t_R port map( A => crossbar_in(132), Y => n858);
   U1307 : INVx1_ASAP7_75t_R port map( A => crossbar_in(131), Y => n859);
   U1308 : INVx1_ASAP7_75t_R port map( A => crossbar_in(130), Y => n860);
   U1309 : INVx1_ASAP7_75t_R port map( A => crossbar_in(129), Y => n861);
   U1310 : INVx1_ASAP7_75t_R port map( A => crossbar_in(128), Y => n862);
   U1311 : INVx1_ASAP7_75t_R port map( A => crossbar_in(191), Y => n863);
   U1312 : INVx1_ASAP7_75t_R port map( A => crossbar_in(190), Y => n864);
   U1313 : INVx1_ASAP7_75t_R port map( A => crossbar_in(189), Y => n865);
   U1314 : INVx1_ASAP7_75t_R port map( A => crossbar_in(188), Y => n866);
   U1315 : INVx1_ASAP7_75t_R port map( A => crossbar_in(187), Y => n867);
   U1316 : INVx1_ASAP7_75t_R port map( A => crossbar_in(186), Y => n868);
   U1317 : INVx1_ASAP7_75t_R port map( A => crossbar_in(185), Y => n869);
   U1318 : INVx1_ASAP7_75t_R port map( A => crossbar_in(184), Y => n870);
   U1319 : INVx1_ASAP7_75t_R port map( A => crossbar_in(183), Y => n871);
   U1320 : INVx1_ASAP7_75t_R port map( A => crossbar_in(182), Y => n872);
   U1321 : INVx1_ASAP7_75t_R port map( A => crossbar_in(181), Y => n873);
   U1322 : INVx1_ASAP7_75t_R port map( A => crossbar_in(180), Y => n874);
   U1323 : INVx1_ASAP7_75t_R port map( A => crossbar_in(179), Y => n875);
   U1324 : INVx1_ASAP7_75t_R port map( A => crossbar_in(178), Y => n876);
   U1325 : INVx1_ASAP7_75t_R port map( A => crossbar_in(177), Y => n877);
   U1326 : INVx1_ASAP7_75t_R port map( A => crossbar_in(176), Y => n878);
   U1327 : INVx1_ASAP7_75t_R port map( A => crossbar_in(175), Y => n879);
   U1328 : INVx1_ASAP7_75t_R port map( A => crossbar_in(174), Y => n880);
   U1329 : INVx1_ASAP7_75t_R port map( A => crossbar_in(173), Y => n881);
   U1330 : INVx1_ASAP7_75t_R port map( A => crossbar_in(172), Y => n882);
   U1331 : INVx1_ASAP7_75t_R port map( A => crossbar_in(171), Y => n883);
   U1332 : INVx1_ASAP7_75t_R port map( A => crossbar_in(170), Y => n884);
   U1333 : INVx1_ASAP7_75t_R port map( A => crossbar_in(169), Y => n885);
   U1334 : INVx1_ASAP7_75t_R port map( A => crossbar_in(168), Y => n886);
   U1335 : INVx1_ASAP7_75t_R port map( A => crossbar_in(167), Y => n887);
   U1336 : INVx1_ASAP7_75t_R port map( A => crossbar_in(166), Y => n888);
   U1337 : INVx1_ASAP7_75t_R port map( A => crossbar_in(165), Y => n889);
   U1338 : INVx1_ASAP7_75t_R port map( A => crossbar_in(164), Y => n890);
   U1339 : INVx1_ASAP7_75t_R port map( A => crossbar_in(163), Y => n891);
   U1340 : INVx1_ASAP7_75t_R port map( A => crossbar_in(162), Y => n892);
   U1341 : INVx1_ASAP7_75t_R port map( A => crossbar_in(161), Y => n893);
   U1342 : INVx1_ASAP7_75t_R port map( A => crossbar_in(160), Y => n894);
   U1343 : INVx1_ASAP7_75t_R port map( A => crossbar_in(159), Y => n895);
   U1344 : INVx1_ASAP7_75t_R port map( A => crossbar_in(158), Y => n896);
   U1345 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(17), Y => n897);
   U1346 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(16), Y => n898);
   U1347 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(15), Y => n899);
   U1348 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(10), Y => n900);
   U1349 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(11), Y => n901);
   U1350 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(9), Y => n902);
   U1351 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(14), Y => n903);
   U1352 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(13), Y => n904);
   U1353 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(5), Y => n905);
   U1354 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(4), Y => n906);
   U1355 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(3), Y => n907);
   U1356 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(7), Y => n908);
   U1357 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(8), Y => n909);
   U1358 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(6), Y => n910);
   U1359 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(2), Y => n911);
   U1360 : INVx1_ASAP7_75t_R port map( A => crossbar_ctrl(1), Y => n912);
   U1361 : INVx1_ASAP7_75t_R port map( A => crossbar_in(0), Y => n913);
   U1362 : INVx1_ASAP7_75t_R port map( A => crossbar_in(10), Y => n914);
   U1363 : INVx1_ASAP7_75t_R port map( A => crossbar_in(11), Y => n915);
   U1364 : INVx1_ASAP7_75t_R port map( A => crossbar_in(12), Y => n916);
   U1365 : INVx1_ASAP7_75t_R port map( A => crossbar_in(13), Y => n917);
   U1366 : INVx1_ASAP7_75t_R port map( A => crossbar_in(14), Y => n918);
   U1367 : INVx1_ASAP7_75t_R port map( A => crossbar_in(15), Y => n919);
   U1368 : INVx1_ASAP7_75t_R port map( A => crossbar_in(16), Y => n920);
   U1369 : INVx1_ASAP7_75t_R port map( A => crossbar_in(17), Y => n921);
   U1370 : INVx1_ASAP7_75t_R port map( A => crossbar_in(18), Y => n922);
   U1371 : INVx1_ASAP7_75t_R port map( A => crossbar_in(19), Y => n923);
   U1372 : INVx1_ASAP7_75t_R port map( A => crossbar_in(1), Y => n924);
   U1373 : INVx1_ASAP7_75t_R port map( A => crossbar_in(20), Y => n925);
   U1374 : INVx1_ASAP7_75t_R port map( A => crossbar_in(21), Y => n926);
   U1375 : INVx1_ASAP7_75t_R port map( A => crossbar_in(22), Y => n927);
   U1376 : INVx1_ASAP7_75t_R port map( A => crossbar_in(23), Y => n928);
   U1377 : INVx1_ASAP7_75t_R port map( A => crossbar_in(24), Y => n929);
   U1378 : INVx1_ASAP7_75t_R port map( A => crossbar_in(25), Y => n930);
   U1379 : INVx1_ASAP7_75t_R port map( A => crossbar_in(26), Y => n931);
   U1380 : INVx1_ASAP7_75t_R port map( A => crossbar_in(27), Y => n932);
   U1381 : INVx1_ASAP7_75t_R port map( A => crossbar_in(28), Y => n933);
   U1382 : INVx1_ASAP7_75t_R port map( A => crossbar_in(29), Y => n934);
   U1383 : INVx1_ASAP7_75t_R port map( A => crossbar_in(2), Y => n935);
   U1384 : INVx1_ASAP7_75t_R port map( A => crossbar_in(30), Y => n936);
   U1385 : INVx1_ASAP7_75t_R port map( A => crossbar_in(31), Y => n937);
   U1386 : INVx1_ASAP7_75t_R port map( A => crossbar_in(32), Y => n938);
   U1387 : INVx1_ASAP7_75t_R port map( A => crossbar_in(33), Y => n939);
   U1388 : INVx1_ASAP7_75t_R port map( A => crossbar_in(34), Y => n940);
   U1389 : INVx1_ASAP7_75t_R port map( A => crossbar_in(35), Y => n941);
   U1390 : INVx1_ASAP7_75t_R port map( A => crossbar_in(36), Y => n942);
   U1391 : INVx1_ASAP7_75t_R port map( A => crossbar_in(37), Y => n943);
   U1392 : INVx1_ASAP7_75t_R port map( A => crossbar_in(38), Y => n944);
   U1393 : INVx1_ASAP7_75t_R port map( A => crossbar_in(39), Y => n945);
   U1394 : INVx1_ASAP7_75t_R port map( A => crossbar_in(3), Y => n946);
   U1395 : INVx1_ASAP7_75t_R port map( A => crossbar_in(40), Y => n947);
   U1396 : INVx1_ASAP7_75t_R port map( A => crossbar_in(41), Y => n948);
   U1397 : INVx1_ASAP7_75t_R port map( A => crossbar_in(42), Y => n949);
   U1398 : INVx1_ASAP7_75t_R port map( A => crossbar_in(43), Y => n950);
   U1399 : INVx1_ASAP7_75t_R port map( A => crossbar_in(44), Y => n951);
   U1400 : INVx1_ASAP7_75t_R port map( A => crossbar_in(45), Y => n952);
   U1401 : INVx1_ASAP7_75t_R port map( A => crossbar_in(46), Y => n953);
   U1402 : INVx1_ASAP7_75t_R port map( A => crossbar_in(47), Y => n954);
   U1403 : INVx1_ASAP7_75t_R port map( A => crossbar_in(48), Y => n955);
   U1404 : INVx1_ASAP7_75t_R port map( A => crossbar_in(49), Y => n956);
   U1405 : INVx1_ASAP7_75t_R port map( A => crossbar_in(4), Y => n957);
   U1406 : INVx1_ASAP7_75t_R port map( A => crossbar_in(50), Y => n958);
   U1407 : INVx1_ASAP7_75t_R port map( A => crossbar_in(51), Y => n959);
   U1408 : INVx1_ASAP7_75t_R port map( A => crossbar_in(52), Y => n960);
   U1409 : INVx1_ASAP7_75t_R port map( A => crossbar_in(53), Y => n961);
   U1410 : INVx1_ASAP7_75t_R port map( A => crossbar_in(54), Y => n962);
   U1411 : INVx1_ASAP7_75t_R port map( A => crossbar_in(55), Y => n963);
   U1412 : INVx1_ASAP7_75t_R port map( A => crossbar_in(56), Y => n964);
   U1413 : INVx1_ASAP7_75t_R port map( A => crossbar_in(57), Y => n965);
   U1414 : INVx1_ASAP7_75t_R port map( A => crossbar_in(58), Y => n966);
   U1415 : INVx1_ASAP7_75t_R port map( A => crossbar_in(59), Y => n967);
   U1416 : INVx1_ASAP7_75t_R port map( A => crossbar_in(5), Y => n968);
   U1417 : INVx1_ASAP7_75t_R port map( A => crossbar_in(60), Y => n969);
   U1418 : INVx1_ASAP7_75t_R port map( A => crossbar_in(61), Y => n970);
   U1419 : INVx1_ASAP7_75t_R port map( A => crossbar_in(62), Y => n971);
   U1420 : INVx1_ASAP7_75t_R port map( A => crossbar_in(63), Y => n972);
   U1421 : INVx1_ASAP7_75t_R port map( A => crossbar_in(6), Y => n973);
   U1422 : INVx1_ASAP7_75t_R port map( A => crossbar_in(7), Y => n974);
   U1423 : INVx1_ASAP7_75t_R port map( A => crossbar_in(8), Y => n975);
   U1424 : INVx1_ASAP7_75t_R port map( A => crossbar_in(9), Y => n976);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity vc_input_buffer_2_0000000200000002_0 is

   port( clk, rst : in std_logic;  data_rx : in std_logic_vector (63 downto 0);
         vc_write_rx, vc_transfer : in std_logic_vector (1 downto 0);  
         valid_data_vc : out std_logic_vector (1 downto 0);  data_transfer : 
         out std_logic_vector (63 downto 0);  header : out std_logic_vector (19
         downto 0));

end vc_input_buffer_2_0000000200000002_0;

architecture SYN_rtl of vc_input_buffer_2_0000000200000002_0 is

   component HB1xp67_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVx1_ASAP7_75t_R
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component fifo_buff_depth2_11
      port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, 
            clk, rst : in std_logic;  data_out : out std_logic_vector (63 
            downto 0);  valid_data : out std_logic);
   end component;
   
   component fifo_buff_depth2_12
      port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, 
            clk, rst : in std_logic;  data_out : out std_logic_vector (63 
            downto 0);  valid_data : out std_logic);
   end component;
   
   component AO22x1_ASAP7_75t_R
      port( A1, A2, B1, B2 : in std_logic;  Y : out std_logic);
   end component;
   
   signal header_1_PACKET_LENGTH_3_port, header_1_PACKET_LENGTH_2_port, 
      header_1_PACKET_LENGTH_1_port, header_1_PACKET_LENGTH_0_port, 
      header_1_X_DEST_1_port, header_1_X_DEST_0_port, header_1_Y_DEST_1_port, 
      header_1_Y_DEST_0_port, header_1_Z_DEST_1_port, header_1_Z_DEST_0_port, 
      header_0_PACKET_LENGTH_3_port, header_0_PACKET_LENGTH_2_port, 
      header_0_PACKET_LENGTH_1_port, header_0_PACKET_LENGTH_0_port, 
      header_0_X_DEST_1_port, header_0_X_DEST_0_port, header_0_Y_DEST_1_port, 
      header_0_Y_DEST_0_port, header_0_Z_DEST_1_port, header_0_Z_DEST_0_port, 
      buffer_out_vector_1_63_port, buffer_out_vector_1_62_port, 
      buffer_out_vector_1_61_port, buffer_out_vector_1_60_port, 
      buffer_out_vector_1_59_port, buffer_out_vector_1_58_port, 
      buffer_out_vector_1_57_port, buffer_out_vector_1_56_port, 
      buffer_out_vector_1_55_port, buffer_out_vector_1_54_port, 
      buffer_out_vector_1_53_port, buffer_out_vector_1_52_port, 
      buffer_out_vector_1_51_port, buffer_out_vector_1_50_port, 
      buffer_out_vector_1_49_port, buffer_out_vector_1_48_port, 
      buffer_out_vector_1_47_port, buffer_out_vector_1_46_port, 
      buffer_out_vector_1_45_port, buffer_out_vector_1_44_port, 
      buffer_out_vector_1_43_port, buffer_out_vector_1_42_port, 
      buffer_out_vector_1_41_port, buffer_out_vector_1_40_port, 
      buffer_out_vector_1_39_port, buffer_out_vector_1_38_port, 
      buffer_out_vector_1_37_port, buffer_out_vector_1_36_port, 
      buffer_out_vector_1_35_port, buffer_out_vector_1_34_port, 
      buffer_out_vector_1_33_port, buffer_out_vector_1_32_port, 
      buffer_out_vector_1_31_port, buffer_out_vector_1_30_port, 
      buffer_out_vector_1_29_port, buffer_out_vector_1_28_port, 
      buffer_out_vector_1_27_port, buffer_out_vector_1_26_port, 
      buffer_out_vector_1_25_port, buffer_out_vector_1_24_port, 
      buffer_out_vector_1_23_port, buffer_out_vector_1_22_port, 
      buffer_out_vector_1_21_port, buffer_out_vector_1_20_port, 
      buffer_out_vector_1_19_port, buffer_out_vector_1_18_port, 
      buffer_out_vector_1_17_port, buffer_out_vector_1_16_port, 
      buffer_out_vector_1_15_port, buffer_out_vector_1_14_port, 
      buffer_out_vector_1_13_port, buffer_out_vector_1_12_port, 
      buffer_out_vector_1_11_port, buffer_out_vector_1_10_port, 
      buffer_out_vector_0_63_port, buffer_out_vector_0_62_port, 
      buffer_out_vector_0_61_port, buffer_out_vector_0_60_port, 
      buffer_out_vector_0_59_port, buffer_out_vector_0_58_port, 
      buffer_out_vector_0_57_port, buffer_out_vector_0_56_port, 
      buffer_out_vector_0_55_port, buffer_out_vector_0_54_port, 
      buffer_out_vector_0_53_port, buffer_out_vector_0_52_port, 
      buffer_out_vector_0_51_port, buffer_out_vector_0_50_port, 
      buffer_out_vector_0_49_port, buffer_out_vector_0_48_port, 
      buffer_out_vector_0_47_port, buffer_out_vector_0_46_port, 
      buffer_out_vector_0_45_port, buffer_out_vector_0_44_port, 
      buffer_out_vector_0_43_port, buffer_out_vector_0_42_port, 
      buffer_out_vector_0_41_port, buffer_out_vector_0_40_port, 
      buffer_out_vector_0_39_port, buffer_out_vector_0_38_port, 
      buffer_out_vector_0_37_port, buffer_out_vector_0_36_port, 
      buffer_out_vector_0_35_port, buffer_out_vector_0_34_port, 
      buffer_out_vector_0_33_port, buffer_out_vector_0_32_port, 
      buffer_out_vector_0_31_port, buffer_out_vector_0_30_port, 
      buffer_out_vector_0_29_port, buffer_out_vector_0_28_port, 
      buffer_out_vector_0_27_port, buffer_out_vector_0_26_port, 
      buffer_out_vector_0_25_port, buffer_out_vector_0_24_port, 
      buffer_out_vector_0_23_port, buffer_out_vector_0_22_port, 
      buffer_out_vector_0_21_port, buffer_out_vector_0_20_port, 
      buffer_out_vector_0_19_port, buffer_out_vector_0_18_port, 
      buffer_out_vector_0_17_port, buffer_out_vector_0_16_port, 
      buffer_out_vector_0_15_port, buffer_out_vector_0_14_port, 
      buffer_out_vector_0_13_port, buffer_out_vector_0_12_port, 
      buffer_out_vector_0_11_port, buffer_out_vector_0_10_port, n1, n2, n3, n4,
      n5, n6, n7, n8 : std_logic;

begin
   header <= ( header_1_PACKET_LENGTH_3_port, header_1_PACKET_LENGTH_2_port, 
      header_1_PACKET_LENGTH_1_port, header_1_PACKET_LENGTH_0_port, 
      header_1_X_DEST_1_port, header_1_X_DEST_0_port, header_1_Y_DEST_1_port, 
      header_1_Y_DEST_0_port, header_1_Z_DEST_1_port, header_1_Z_DEST_0_port, 
      header_0_PACKET_LENGTH_3_port, header_0_PACKET_LENGTH_2_port, 
      header_0_PACKET_LENGTH_1_port, header_0_PACKET_LENGTH_0_port, 
      header_0_X_DEST_1_port, header_0_X_DEST_0_port, header_0_Y_DEST_1_port, 
      header_0_Y_DEST_0_port, header_0_Z_DEST_1_port, header_0_Z_DEST_0_port );
   
   U2 : AO22x1_ASAP7_75t_R port map( A1 => n3, A2 => 
                           buffer_out_vector_1_30_port, B1 => 
                           buffer_out_vector_0_30_port, B2 => n4, Y => 
                           data_transfer(30));
   U3 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_31_port, A2 => 
                           n3, B1 => buffer_out_vector_0_31_port, B2 => n4, Y 
                           => data_transfer(31));
   U4 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_32_port, A2 => 
                           n3, B1 => buffer_out_vector_0_32_port, B2 => n4, Y 
                           => data_transfer(32));
   U5 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_33_port, A2 => 
                           n3, B1 => buffer_out_vector_0_33_port, B2 => n4, Y 
                           => data_transfer(33));
   U6 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_34_port, A2 => 
                           n3, B1 => buffer_out_vector_0_34_port, B2 => n4, Y 
                           => data_transfer(34));
   U7 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_35_port, A2 => 
                           n3, B1 => buffer_out_vector_0_35_port, B2 => n6, Y 
                           => data_transfer(35));
   U8 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_36_port, A2 => 
                           n3, B1 => buffer_out_vector_0_36_port, B2 => n5, Y 
                           => data_transfer(36));
   U9 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_37_port, A2 => 
                           n3, B1 => buffer_out_vector_0_37_port, B2 => n7, Y 
                           => data_transfer(37));
   U10 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_38_port, A2 => 
                           n3, B1 => buffer_out_vector_0_38_port, B2 => n6, Y 
                           => data_transfer(38));
   U11 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_39_port, A2 => 
                           n3, B1 => buffer_out_vector_0_39_port, B2 => n5, Y 
                           => data_transfer(39));
   U12 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_40_port, A2 => 
                           n3, B1 => buffer_out_vector_0_40_port, B2 => n7, Y 
                           => data_transfer(40));
   U13 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_41_port, A2 => 
                           n3, B1 => buffer_out_vector_0_41_port, B2 => n6, Y 
                           => data_transfer(41));
   U14 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_42_port, A2 => 
                           n3, B1 => buffer_out_vector_0_42_port, B2 => n5, Y 
                           => data_transfer(42));
   U15 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_43_port, A2 => 
                           n3, B1 => buffer_out_vector_0_43_port, B2 => n7, Y 
                           => data_transfer(43));
   U16 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_44_port, A2 => 
                           n3, B1 => buffer_out_vector_0_44_port, B2 => n7, Y 
                           => data_transfer(44));
   U17 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_45_port, A2 => 
                           n3, B1 => buffer_out_vector_0_45_port, B2 => n6, Y 
                           => data_transfer(45));
   U18 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_46_port, A2 => 
                           n3, B1 => buffer_out_vector_0_46_port, B2 => n5, Y 
                           => data_transfer(46));
   U19 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_47_port, A2 => 
                           n3, B1 => buffer_out_vector_0_47_port, B2 => n6, Y 
                           => data_transfer(47));
   U20 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_48_port, A2 => 
                           n3, B1 => buffer_out_vector_0_48_port, B2 => n6, Y 
                           => data_transfer(48));
   U21 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_49_port, A2 => 
                           n3, B1 => buffer_out_vector_0_49_port, B2 => n7, Y 
                           => data_transfer(49));
   U22 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_50_port, A2 => 
                           n3, B1 => buffer_out_vector_0_50_port, B2 => n6, Y 
                           => data_transfer(50));
   U23 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_51_port, A2 => 
                           n2, B1 => buffer_out_vector_0_51_port, B2 => n7, Y 
                           => data_transfer(51));
   U24 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_52_port, A2 => 
                           n2, B1 => buffer_out_vector_0_52_port, B2 => n5, Y 
                           => data_transfer(52));
   U25 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_53_port, A2 => 
                           n2, B1 => buffer_out_vector_0_53_port, B2 => n6, Y 
                           => data_transfer(53));
   U26 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_54_port, A2 => 
                           n2, B1 => buffer_out_vector_0_54_port, B2 => n7, Y 
                           => data_transfer(54));
   U27 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_55_port, A2 => 
                           n2, B1 => buffer_out_vector_0_55_port, B2 => n6, Y 
                           => data_transfer(55));
   U28 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_56_port, A2 => 
                           n2, B1 => buffer_out_vector_0_56_port, B2 => n5, Y 
                           => data_transfer(56));
   U29 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_57_port, A2 => 
                           n2, B1 => buffer_out_vector_0_57_port, B2 => n7, Y 
                           => data_transfer(57));
   U30 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_58_port, A2 => 
                           n2, B1 => buffer_out_vector_0_58_port, B2 => n6, Y 
                           => data_transfer(58));
   U31 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_59_port, A2 => 
                           n2, B1 => buffer_out_vector_0_59_port, B2 => n5, Y 
                           => data_transfer(59));
   U32 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_60_port, A2 => 
                           n2, B1 => buffer_out_vector_0_60_port, B2 => n6, Y 
                           => data_transfer(60));
   U33 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_61_port, A2 => 
                           n2, B1 => buffer_out_vector_0_61_port, B2 => n7, Y 
                           => data_transfer(61));
   U34 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_62_port, A2 => 
                           n2, B1 => buffer_out_vector_0_62_port, B2 => n6, Y 
                           => data_transfer(62));
   U35 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_63_port, A2 => 
                           n2, B1 => buffer_out_vector_0_63_port, B2 => n5, Y 
                           => data_transfer(63));
   U36 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_0_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_0_port, B2 => n7
                           , Y => data_transfer(0));
   U37 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_1_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_1_port, B2 => n5
                           , Y => data_transfer(1));
   U38 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_2_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_2_port, B2 => n7
                           , Y => data_transfer(2));
   U39 : AO22x1_ASAP7_75t_R port map( A1 => header_1_PACKET_LENGTH_3_port, A2 
                           => n2, B1 => header_0_PACKET_LENGTH_3_port, B2 => n5
                           , Y => data_transfer(3));
   U40 : AO22x1_ASAP7_75t_R port map( A1 => header_1_X_DEST_0_port, A2 => n2, 
                           B1 => header_0_X_DEST_0_port, B2 => n5, Y => 
                           data_transfer(4));
   U41 : AO22x1_ASAP7_75t_R port map( A1 => header_1_X_DEST_1_port, A2 => n2, 
                           B1 => header_0_X_DEST_1_port, B2 => n5, Y => 
                           data_transfer(5));
   U42 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Y_DEST_0_port, A2 => n2, 
                           B1 => header_0_Y_DEST_0_port, B2 => n5, Y => 
                           data_transfer(6));
   U43 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Y_DEST_1_port, A2 => n2, 
                           B1 => header_0_Y_DEST_1_port, B2 => n5, Y => 
                           data_transfer(7));
   U44 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Z_DEST_0_port, A2 => n2, 
                           B1 => header_0_Z_DEST_0_port, B2 => n5, Y => 
                           data_transfer(8));
   U45 : AO22x1_ASAP7_75t_R port map( A1 => header_1_Z_DEST_1_port, A2 => n2, 
                           B1 => header_0_Z_DEST_1_port, B2 => n5, Y => 
                           data_transfer(9));
   U46 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_10_port, A2 => 
                           n2, B1 => buffer_out_vector_0_10_port, B2 => n5, Y 
                           => data_transfer(10));
   U47 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_11_port, A2 => 
                           n2, B1 => buffer_out_vector_0_11_port, B2 => n6, Y 
                           => data_transfer(11));
   U48 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_12_port, A2 => 
                           n2, B1 => buffer_out_vector_0_12_port, B2 => n6, Y 
                           => data_transfer(12));
   U49 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_13_port, A2 => 
                           n2, B1 => buffer_out_vector_0_13_port, B2 => n6, Y 
                           => data_transfer(13));
   U50 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_14_port, A2 => 
                           n2, B1 => buffer_out_vector_0_14_port, B2 => n6, Y 
                           => data_transfer(14));
   U51 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_15_port, A2 => 
                           n2, B1 => buffer_out_vector_0_15_port, B2 => n6, Y 
                           => data_transfer(15));
   U52 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_16_port, A2 => 
                           n2, B1 => buffer_out_vector_0_16_port, B2 => n6, Y 
                           => data_transfer(16));
   U53 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_17_port, A2 => 
                           n2, B1 => buffer_out_vector_0_17_port, B2 => n6, Y 
                           => data_transfer(17));
   U54 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_18_port, A2 => 
                           n2, B1 => buffer_out_vector_0_18_port, B2 => n6, Y 
                           => data_transfer(18));
   U55 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_19_port, A2 => 
                           n2, B1 => buffer_out_vector_0_19_port, B2 => n7, Y 
                           => data_transfer(19));
   U56 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_20_port, A2 => 
                           n2, B1 => buffer_out_vector_0_20_port, B2 => n7, Y 
                           => data_transfer(20));
   U57 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_21_port, A2 => 
                           n2, B1 => buffer_out_vector_0_21_port, B2 => n7, Y 
                           => data_transfer(21));
   U58 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_22_port, A2 => 
                           n2, B1 => buffer_out_vector_0_22_port, B2 => n7, Y 
                           => data_transfer(22));
   U59 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_23_port, A2 => 
                           n2, B1 => buffer_out_vector_0_23_port, B2 => n7, Y 
                           => data_transfer(23));
   U60 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_24_port, A2 => 
                           n2, B1 => buffer_out_vector_0_24_port, B2 => n7, Y 
                           => data_transfer(24));
   U61 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_25_port, A2 => 
                           n2, B1 => buffer_out_vector_0_25_port, B2 => n7, Y 
                           => data_transfer(25));
   U62 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_26_port, A2 => 
                           n2, B1 => buffer_out_vector_0_26_port, B2 => n7, Y 
                           => data_transfer(26));
   U63 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_27_port, A2 => 
                           n2, B1 => buffer_out_vector_0_27_port, B2 => n5, Y 
                           => data_transfer(27));
   U64 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_28_port, A2 => 
                           n2, B1 => buffer_out_vector_0_28_port, B2 => n5, Y 
                           => data_transfer(28));
   U65 : AO22x1_ASAP7_75t_R port map( A1 => buffer_out_vector_1_29_port, A2 => 
                           n2, B1 => buffer_out_vector_0_29_port, B2 => n5, Y 
                           => data_transfer(29));
   fifo_i_0 : fifo_buff_depth2_12 port map( data_in(63) => data_rx(63), 
                           data_in(62) => data_rx(62), data_in(61) => 
                           data_rx(61), data_in(60) => data_rx(60), data_in(59)
                           => data_rx(59), data_in(58) => data_rx(58), 
                           data_in(57) => data_rx(57), data_in(56) => 
                           data_rx(56), data_in(55) => data_rx(55), data_in(54)
                           => data_rx(54), data_in(53) => data_rx(53), 
                           data_in(52) => data_rx(52), data_in(51) => 
                           data_rx(51), data_in(50) => data_rx(50), data_in(49)
                           => data_rx(49), data_in(48) => data_rx(48), 
                           data_in(47) => data_rx(47), data_in(46) => 
                           data_rx(46), data_in(45) => data_rx(45), data_in(44)
                           => data_rx(44), data_in(43) => data_rx(43), 
                           data_in(42) => data_rx(42), data_in(41) => 
                           data_rx(41), data_in(40) => data_rx(40), data_in(39)
                           => data_rx(39), data_in(38) => data_rx(38), 
                           data_in(37) => data_rx(37), data_in(36) => 
                           data_rx(36), data_in(35) => data_rx(35), data_in(34)
                           => data_rx(34), data_in(33) => data_rx(33), 
                           data_in(32) => data_rx(32), data_in(31) => 
                           data_rx(31), data_in(30) => data_rx(30), data_in(29)
                           => data_rx(29), data_in(28) => data_rx(28), 
                           data_in(27) => data_rx(27), data_in(26) => 
                           data_rx(26), data_in(25) => data_rx(25), data_in(24)
                           => data_rx(24), data_in(23) => data_rx(23), 
                           data_in(22) => data_rx(22), data_in(21) => 
                           data_rx(21), data_in(20) => data_rx(20), data_in(19)
                           => data_rx(19), data_in(18) => data_rx(18), 
                           data_in(17) => data_rx(17), data_in(16) => 
                           data_rx(16), data_in(15) => data_rx(15), data_in(14)
                           => data_rx(14), data_in(13) => data_rx(13), 
                           data_in(12) => data_rx(12), data_in(11) => 
                           data_rx(11), data_in(10) => data_rx(10), data_in(9) 
                           => data_rx(9), data_in(8) => data_rx(8), data_in(7) 
                           => data_rx(7), data_in(6) => data_rx(6), data_in(5) 
                           => data_rx(5), data_in(4) => data_rx(4), data_in(3) 
                           => data_rx(3), data_in(2) => data_rx(2), data_in(1) 
                           => data_rx(1), data_in(0) => data_rx(0), write_en =>
                           vc_write_rx(0), read_en => vc_transfer(0), clk => 
                           clk, rst => n8, data_out(63) => 
                           buffer_out_vector_0_63_port, data_out(62) => 
                           buffer_out_vector_0_62_port, data_out(61) => 
                           buffer_out_vector_0_61_port, data_out(60) => 
                           buffer_out_vector_0_60_port, data_out(59) => 
                           buffer_out_vector_0_59_port, data_out(58) => 
                           buffer_out_vector_0_58_port, data_out(57) => 
                           buffer_out_vector_0_57_port, data_out(56) => 
                           buffer_out_vector_0_56_port, data_out(55) => 
                           buffer_out_vector_0_55_port, data_out(54) => 
                           buffer_out_vector_0_54_port, data_out(53) => 
                           buffer_out_vector_0_53_port, data_out(52) => 
                           buffer_out_vector_0_52_port, data_out(51) => 
                           buffer_out_vector_0_51_port, data_out(50) => 
                           buffer_out_vector_0_50_port, data_out(49) => 
                           buffer_out_vector_0_49_port, data_out(48) => 
                           buffer_out_vector_0_48_port, data_out(47) => 
                           buffer_out_vector_0_47_port, data_out(46) => 
                           buffer_out_vector_0_46_port, data_out(45) => 
                           buffer_out_vector_0_45_port, data_out(44) => 
                           buffer_out_vector_0_44_port, data_out(43) => 
                           buffer_out_vector_0_43_port, data_out(42) => 
                           buffer_out_vector_0_42_port, data_out(41) => 
                           buffer_out_vector_0_41_port, data_out(40) => 
                           buffer_out_vector_0_40_port, data_out(39) => 
                           buffer_out_vector_0_39_port, data_out(38) => 
                           buffer_out_vector_0_38_port, data_out(37) => 
                           buffer_out_vector_0_37_port, data_out(36) => 
                           buffer_out_vector_0_36_port, data_out(35) => 
                           buffer_out_vector_0_35_port, data_out(34) => 
                           buffer_out_vector_0_34_port, data_out(33) => 
                           buffer_out_vector_0_33_port, data_out(32) => 
                           buffer_out_vector_0_32_port, data_out(31) => 
                           buffer_out_vector_0_31_port, data_out(30) => 
                           buffer_out_vector_0_30_port, data_out(29) => 
                           buffer_out_vector_0_29_port, data_out(28) => 
                           buffer_out_vector_0_28_port, data_out(27) => 
                           buffer_out_vector_0_27_port, data_out(26) => 
                           buffer_out_vector_0_26_port, data_out(25) => 
                           buffer_out_vector_0_25_port, data_out(24) => 
                           buffer_out_vector_0_24_port, data_out(23) => 
                           buffer_out_vector_0_23_port, data_out(22) => 
                           buffer_out_vector_0_22_port, data_out(21) => 
                           buffer_out_vector_0_21_port, data_out(20) => 
                           buffer_out_vector_0_20_port, data_out(19) => 
                           buffer_out_vector_0_19_port, data_out(18) => 
                           buffer_out_vector_0_18_port, data_out(17) => 
                           buffer_out_vector_0_17_port, data_out(16) => 
                           buffer_out_vector_0_16_port, data_out(15) => 
                           buffer_out_vector_0_15_port, data_out(14) => 
                           buffer_out_vector_0_14_port, data_out(13) => 
                           buffer_out_vector_0_13_port, data_out(12) => 
                           buffer_out_vector_0_12_port, data_out(11) => 
                           buffer_out_vector_0_11_port, data_out(10) => 
                           buffer_out_vector_0_10_port, data_out(9) => 
                           header_0_Z_DEST_1_port, data_out(8) => 
                           header_0_Z_DEST_0_port, data_out(7) => 
                           header_0_Y_DEST_1_port, data_out(6) => 
                           header_0_Y_DEST_0_port, data_out(5) => 
                           header_0_X_DEST_1_port, data_out(4) => 
                           header_0_X_DEST_0_port, data_out(3) => 
                           header_0_PACKET_LENGTH_3_port, data_out(2) => 
                           header_0_PACKET_LENGTH_2_port, data_out(1) => 
                           header_0_PACKET_LENGTH_1_port, data_out(0) => 
                           header_0_PACKET_LENGTH_0_port, valid_data => 
                           valid_data_vc(0));
   fifo_i_1 : fifo_buff_depth2_11 port map( data_in(63) => data_rx(63), 
                           data_in(62) => data_rx(62), data_in(61) => 
                           data_rx(61), data_in(60) => data_rx(60), data_in(59)
                           => data_rx(59), data_in(58) => data_rx(58), 
                           data_in(57) => data_rx(57), data_in(56) => 
                           data_rx(56), data_in(55) => data_rx(55), data_in(54)
                           => data_rx(54), data_in(53) => data_rx(53), 
                           data_in(52) => data_rx(52), data_in(51) => 
                           data_rx(51), data_in(50) => data_rx(50), data_in(49)
                           => data_rx(49), data_in(48) => data_rx(48), 
                           data_in(47) => data_rx(47), data_in(46) => 
                           data_rx(46), data_in(45) => data_rx(45), data_in(44)
                           => data_rx(44), data_in(43) => data_rx(43), 
                           data_in(42) => data_rx(42), data_in(41) => 
                           data_rx(41), data_in(40) => data_rx(40), data_in(39)
                           => data_rx(39), data_in(38) => data_rx(38), 
                           data_in(37) => data_rx(37), data_in(36) => 
                           data_rx(36), data_in(35) => data_rx(35), data_in(34)
                           => data_rx(34), data_in(33) => data_rx(33), 
                           data_in(32) => data_rx(32), data_in(31) => 
                           data_rx(31), data_in(30) => data_rx(30), data_in(29)
                           => data_rx(29), data_in(28) => data_rx(28), 
                           data_in(27) => data_rx(27), data_in(26) => 
                           data_rx(26), data_in(25) => data_rx(25), data_in(24)
                           => data_rx(24), data_in(23) => data_rx(23), 
                           data_in(22) => data_rx(22), data_in(21) => 
                           data_rx(21), data_in(20) => data_rx(20), data_in(19)
                           => data_rx(19), data_in(18) => data_rx(18), 
                           data_in(17) => data_rx(17), data_in(16) => 
                           data_rx(16), data_in(15) => data_rx(15), data_in(14)
                           => data_rx(14), data_in(13) => data_rx(13), 
                           data_in(12) => data_rx(12), data_in(11) => 
                           data_rx(11), data_in(10) => data_rx(10), data_in(9) 
                           => data_rx(9), data_in(8) => data_rx(8), data_in(7) 
                           => data_rx(7), data_in(6) => data_rx(6), data_in(5) 
                           => data_rx(5), data_in(4) => data_rx(4), data_in(3) 
                           => data_rx(3), data_in(2) => data_rx(2), data_in(1) 
                           => data_rx(1), data_in(0) => data_rx(0), write_en =>
                           vc_write_rx(1), read_en => n2, clk => clk, rst => n8
                           , data_out(63) => buffer_out_vector_1_63_port, 
                           data_out(62) => buffer_out_vector_1_62_port, 
                           data_out(61) => buffer_out_vector_1_61_port, 
                           data_out(60) => buffer_out_vector_1_60_port, 
                           data_out(59) => buffer_out_vector_1_59_port, 
                           data_out(58) => buffer_out_vector_1_58_port, 
                           data_out(57) => buffer_out_vector_1_57_port, 
                           data_out(56) => buffer_out_vector_1_56_port, 
                           data_out(55) => buffer_out_vector_1_55_port, 
                           data_out(54) => buffer_out_vector_1_54_port, 
                           data_out(53) => buffer_out_vector_1_53_port, 
                           data_out(52) => buffer_out_vector_1_52_port, 
                           data_out(51) => buffer_out_vector_1_51_port, 
                           data_out(50) => buffer_out_vector_1_50_port, 
                           data_out(49) => buffer_out_vector_1_49_port, 
                           data_out(48) => buffer_out_vector_1_48_port, 
                           data_out(47) => buffer_out_vector_1_47_port, 
                           data_out(46) => buffer_out_vector_1_46_port, 
                           data_out(45) => buffer_out_vector_1_45_port, 
                           data_out(44) => buffer_out_vector_1_44_port, 
                           data_out(43) => buffer_out_vector_1_43_port, 
                           data_out(42) => buffer_out_vector_1_42_port, 
                           data_out(41) => buffer_out_vector_1_41_port, 
                           data_out(40) => buffer_out_vector_1_40_port, 
                           data_out(39) => buffer_out_vector_1_39_port, 
                           data_out(38) => buffer_out_vector_1_38_port, 
                           data_out(37) => buffer_out_vector_1_37_port, 
                           data_out(36) => buffer_out_vector_1_36_port, 
                           data_out(35) => buffer_out_vector_1_35_port, 
                           data_out(34) => buffer_out_vector_1_34_port, 
                           data_out(33) => buffer_out_vector_1_33_port, 
                           data_out(32) => buffer_out_vector_1_32_port, 
                           data_out(31) => buffer_out_vector_1_31_port, 
                           data_out(30) => buffer_out_vector_1_30_port, 
                           data_out(29) => buffer_out_vector_1_29_port, 
                           data_out(28) => buffer_out_vector_1_28_port, 
                           data_out(27) => buffer_out_vector_1_27_port, 
                           data_out(26) => buffer_out_vector_1_26_port, 
                           data_out(25) => buffer_out_vector_1_25_port, 
                           data_out(24) => buffer_out_vector_1_24_port, 
                           data_out(23) => buffer_out_vector_1_23_port, 
                           data_out(22) => buffer_out_vector_1_22_port, 
                           data_out(21) => buffer_out_vector_1_21_port, 
                           data_out(20) => buffer_out_vector_1_20_port, 
                           data_out(19) => buffer_out_vector_1_19_port, 
                           data_out(18) => buffer_out_vector_1_18_port, 
                           data_out(17) => buffer_out_vector_1_17_port, 
                           data_out(16) => buffer_out_vector_1_16_port, 
                           data_out(15) => buffer_out_vector_1_15_port, 
                           data_out(14) => buffer_out_vector_1_14_port, 
                           data_out(13) => buffer_out_vector_1_13_port, 
                           data_out(12) => buffer_out_vector_1_12_port, 
                           data_out(11) => buffer_out_vector_1_11_port, 
                           data_out(10) => buffer_out_vector_1_10_port, 
                           data_out(9) => header_1_Z_DEST_1_port, data_out(8) 
                           => header_1_Z_DEST_0_port, data_out(7) => 
                           header_1_Y_DEST_1_port, data_out(6) => 
                           header_1_Y_DEST_0_port, data_out(5) => 
                           header_1_X_DEST_1_port, data_out(4) => 
                           header_1_X_DEST_0_port, data_out(3) => 
                           header_1_PACKET_LENGTH_3_port, data_out(2) => 
                           header_1_PACKET_LENGTH_2_port, data_out(1) => 
                           header_1_PACKET_LENGTH_1_port, data_out(0) => 
                           header_1_PACKET_LENGTH_0_port, valid_data => 
                           valid_data_vc(1));
   U1 : INVx1_ASAP7_75t_R port map( A => n4, Y => n2);
   U66 : INVx1_ASAP7_75t_R port map( A => n4, Y => n3);
   U67 : INVx1_ASAP7_75t_R port map( A => n1, Y => n4);
   U68 : INVx1_ASAP7_75t_R port map( A => n1, Y => n5);
   U69 : INVx1_ASAP7_75t_R port map( A => n1, Y => n6);
   U70 : INVx1_ASAP7_75t_R port map( A => n1, Y => n7);
   U71 : HB1xp67_ASAP7_75t_R port map( A => vc_transfer(1), Y => n1);
   U72 : HB1xp67_ASAP7_75t_R port map( A => rst, Y => n8);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity vc_input_buffer_1_0000000200000002 is

   port( clk, rst : in std_logic;  data_rx : in std_logic_vector (63 downto 0);
         vc_write_rx, vc_transfer : in std_logic;  valid_data_vc : out 
         std_logic;  data_transfer : out std_logic_vector (63 downto 0);  
         header : out std_logic_vector (9 downto 0));

end vc_input_buffer_1_0000000200000002;

architecture SYN_rtl of vc_input_buffer_1_0000000200000002 is

   component fifo_buff_depth2_0
      port( data_in : in std_logic_vector (63 downto 0);  write_en, read_en, 
            clk, rst : in std_logic;  data_out : out std_logic_vector (63 
            downto 0);  valid_data : out std_logic);
   end component;
   
   signal data_transfer_63_port, data_transfer_62_port, data_transfer_61_port, 
      data_transfer_60_port, data_transfer_59_port, data_transfer_58_port, 
      data_transfer_57_port, data_transfer_56_port, data_transfer_55_port, 
      data_transfer_54_port, data_transfer_53_port, data_transfer_52_port, 
      data_transfer_51_port, data_transfer_50_port, data_transfer_49_port, 
      data_transfer_48_port, data_transfer_47_port, data_transfer_46_port, 
      data_transfer_45_port, data_transfer_44_port, data_transfer_43_port, 
      data_transfer_42_port, data_transfer_41_port, data_transfer_40_port, 
      data_transfer_39_port, data_transfer_38_port, data_transfer_37_port, 
      data_transfer_36_port, data_transfer_35_port, data_transfer_34_port, 
      data_transfer_33_port, data_transfer_32_port, data_transfer_31_port, 
      data_transfer_30_port, data_transfer_29_port, data_transfer_28_port, 
      data_transfer_27_port, data_transfer_26_port, data_transfer_25_port, 
      data_transfer_24_port, data_transfer_23_port, data_transfer_22_port, 
      data_transfer_21_port, data_transfer_20_port, data_transfer_19_port, 
      data_transfer_18_port, data_transfer_17_port, data_transfer_16_port, 
      data_transfer_15_port, data_transfer_14_port, data_transfer_13_port, 
      data_transfer_12_port, data_transfer_11_port, data_transfer_10_port, 
      data_transfer_9_port, data_transfer_8_port, data_transfer_7_port, 
      data_transfer_6_port, data_transfer_5_port, data_transfer_4_port, 
      data_transfer_3_port, data_transfer_2_port, data_transfer_1_port, 
      data_transfer_0_port : std_logic;

begin
   data_transfer <= ( data_transfer_63_port, data_transfer_62_port, 
      data_transfer_61_port, data_transfer_60_port, data_transfer_59_port, 
      data_transfer_58_port, data_transfer_57_port, data_transfer_56_port, 
      data_transfer_55_port, data_transfer_54_port, data_transfer_53_port, 
      data_transfer_52_port, data_transfer_51_port, data_transfer_50_port, 
      data_transfer_49_port, data_transfer_48_port, data_transfer_47_port, 
      data_transfer_46_port, data_transfer_45_port, data_transfer_44_port, 
      data_transfer_43_port, data_transfer_42_port, data_transfer_41_port, 
      data_transfer_40_port, data_transfer_39_port, data_transfer_38_port, 
      data_transfer_37_port, data_transfer_36_port, data_transfer_35_port, 
      data_transfer_34_port, data_transfer_33_port, data_transfer_32_port, 
      data_transfer_31_port, data_transfer_30_port, data_transfer_29_port, 
      data_transfer_28_port, data_transfer_27_port, data_transfer_26_port, 
      data_transfer_25_port, data_transfer_24_port, data_transfer_23_port, 
      data_transfer_22_port, data_transfer_21_port, data_transfer_20_port, 
      data_transfer_19_port, data_transfer_18_port, data_transfer_17_port, 
      data_transfer_16_port, data_transfer_15_port, data_transfer_14_port, 
      data_transfer_13_port, data_transfer_12_port, data_transfer_11_port, 
      data_transfer_10_port, data_transfer_9_port, data_transfer_8_port, 
      data_transfer_7_port, data_transfer_6_port, data_transfer_5_port, 
      data_transfer_4_port, data_transfer_3_port, data_transfer_2_port, 
      data_transfer_1_port, data_transfer_0_port );
   header <= ( data_transfer_3_port, data_transfer_2_port, data_transfer_1_port
      , data_transfer_0_port, data_transfer_5_port, data_transfer_4_port, 
      data_transfer_7_port, data_transfer_6_port, data_transfer_9_port, 
      data_transfer_8_port );
   
   fifo_i_0 : fifo_buff_depth2_0 port map( data_in(63) => data_rx(63), 
                           data_in(62) => data_rx(62), data_in(61) => 
                           data_rx(61), data_in(60) => data_rx(60), data_in(59)
                           => data_rx(59), data_in(58) => data_rx(58), 
                           data_in(57) => data_rx(57), data_in(56) => 
                           data_rx(56), data_in(55) => data_rx(55), data_in(54)
                           => data_rx(54), data_in(53) => data_rx(53), 
                           data_in(52) => data_rx(52), data_in(51) => 
                           data_rx(51), data_in(50) => data_rx(50), data_in(49)
                           => data_rx(49), data_in(48) => data_rx(48), 
                           data_in(47) => data_rx(47), data_in(46) => 
                           data_rx(46), data_in(45) => data_rx(45), data_in(44)
                           => data_rx(44), data_in(43) => data_rx(43), 
                           data_in(42) => data_rx(42), data_in(41) => 
                           data_rx(41), data_in(40) => data_rx(40), data_in(39)
                           => data_rx(39), data_in(38) => data_rx(38), 
                           data_in(37) => data_rx(37), data_in(36) => 
                           data_rx(36), data_in(35) => data_rx(35), data_in(34)
                           => data_rx(34), data_in(33) => data_rx(33), 
                           data_in(32) => data_rx(32), data_in(31) => 
                           data_rx(31), data_in(30) => data_rx(30), data_in(29)
                           => data_rx(29), data_in(28) => data_rx(28), 
                           data_in(27) => data_rx(27), data_in(26) => 
                           data_rx(26), data_in(25) => data_rx(25), data_in(24)
                           => data_rx(24), data_in(23) => data_rx(23), 
                           data_in(22) => data_rx(22), data_in(21) => 
                           data_rx(21), data_in(20) => data_rx(20), data_in(19)
                           => data_rx(19), data_in(18) => data_rx(18), 
                           data_in(17) => data_rx(17), data_in(16) => 
                           data_rx(16), data_in(15) => data_rx(15), data_in(14)
                           => data_rx(14), data_in(13) => data_rx(13), 
                           data_in(12) => data_rx(12), data_in(11) => 
                           data_rx(11), data_in(10) => data_rx(10), data_in(9) 
                           => data_rx(9), data_in(8) => data_rx(8), data_in(7) 
                           => data_rx(7), data_in(6) => data_rx(6), data_in(5) 
                           => data_rx(5), data_in(4) => data_rx(4), data_in(3) 
                           => data_rx(3), data_in(2) => data_rx(2), data_in(1) 
                           => data_rx(1), data_in(0) => data_rx(0), write_en =>
                           vc_write_rx, read_en => vc_transfer, clk => clk, rst
                           => rst, data_out(63) => data_transfer_63_port, 
                           data_out(62) => data_transfer_62_port, data_out(61) 
                           => data_transfer_61_port, data_out(60) => 
                           data_transfer_60_port, data_out(59) => 
                           data_transfer_59_port, data_out(58) => 
                           data_transfer_58_port, data_out(57) => 
                           data_transfer_57_port, data_out(56) => 
                           data_transfer_56_port, data_out(55) => 
                           data_transfer_55_port, data_out(54) => 
                           data_transfer_54_port, data_out(53) => 
                           data_transfer_53_port, data_out(52) => 
                           data_transfer_52_port, data_out(51) => 
                           data_transfer_51_port, data_out(50) => 
                           data_transfer_50_port, data_out(49) => 
                           data_transfer_49_port, data_out(48) => 
                           data_transfer_48_port, data_out(47) => 
                           data_transfer_47_port, data_out(46) => 
                           data_transfer_46_port, data_out(45) => 
                           data_transfer_45_port, data_out(44) => 
                           data_transfer_44_port, data_out(43) => 
                           data_transfer_43_port, data_out(42) => 
                           data_transfer_42_port, data_out(41) => 
                           data_transfer_41_port, data_out(40) => 
                           data_transfer_40_port, data_out(39) => 
                           data_transfer_39_port, data_out(38) => 
                           data_transfer_38_port, data_out(37) => 
                           data_transfer_37_port, data_out(36) => 
                           data_transfer_36_port, data_out(35) => 
                           data_transfer_35_port, data_out(34) => 
                           data_transfer_34_port, data_out(33) => 
                           data_transfer_33_port, data_out(32) => 
                           data_transfer_32_port, data_out(31) => 
                           data_transfer_31_port, data_out(30) => 
                           data_transfer_30_port, data_out(29) => 
                           data_transfer_29_port, data_out(28) => 
                           data_transfer_28_port, data_out(27) => 
                           data_transfer_27_port, data_out(26) => 
                           data_transfer_26_port, data_out(25) => 
                           data_transfer_25_port, data_out(24) => 
                           data_transfer_24_port, data_out(23) => 
                           data_transfer_23_port, data_out(22) => 
                           data_transfer_22_port, data_out(21) => 
                           data_transfer_21_port, data_out(20) => 
                           data_transfer_20_port, data_out(19) => 
                           data_transfer_19_port, data_out(18) => 
                           data_transfer_18_port, data_out(17) => 
                           data_transfer_17_port, data_out(16) => 
                           data_transfer_16_port, data_out(15) => 
                           data_transfer_15_port, data_out(14) => 
                           data_transfer_14_port, data_out(13) => 
                           data_transfer_13_port, data_out(12) => 
                           data_transfer_12_port, data_out(11) => 
                           data_transfer_11_port, data_out(10) => 
                           data_transfer_10_port, data_out(9) => 
                           data_transfer_9_port, data_out(8) => 
                           data_transfer_8_port, data_out(7) => 
                           data_transfer_7_port, data_out(6) => 
                           data_transfer_6_port, data_out(5) => 
                           data_transfer_5_port, data_out(4) => 
                           data_transfer_4_port, data_out(3) => 
                           data_transfer_3_port, data_out(2) => 
                           data_transfer_2_port, data_out(1) => 
                           data_transfer_1_port, data_out(0) => 
                           data_transfer_0_port, valid_data => valid_data_vc);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_router_pl.all;

entity router_pl is

   port( clk, rst : in std_logic;  data_rx : in flit_vector (6 downto 0);  
         vc_write_rx_vec, incr_rx_vec : in std_logic_vector (12 downto 0);  
         data_tx_pl : out flit_vector (6 downto 0);  vc_write_tx_pl_vec, 
         incr_tx_pl_vec : out std_logic_vector (12 downto 0));

end router_pl;

architecture SYN_structural of router_pl is

   component arbiter_7_1_1_1_1_DXYU
      port( clk, rst : in std_logic;  header : in std_logic_vector (129 downto 
            0);  valid_data_vc_vec, incr_rx_vec : in std_logic_vector (12 
            downto 0);  crossbar_ctrl : out std_logic_vector (20 downto 0);  
            vc_transfer_vec, vc_write_tx_vec : out std_logic_vector (12 downto 
            0));
   end component;
   
   component output_register_vc_num2_vc_num_out2_1
      port( clk, rst : in std_logic;  data_tx : in std_logic_vector (63 downto 
            0);  vc_write_tx, incr_tx : in std_logic_vector (1 downto 0);  
            data_tx_pl : out std_logic_vector (63 downto 0);  vc_write_tx_pl, 
            incr_tx_pl : out std_logic_vector (1 downto 0));
   end component;
   
   component output_register_vc_num2_vc_num_out2_2
      port( clk, rst : in std_logic;  data_tx : in std_logic_vector (63 downto 
            0);  vc_write_tx, incr_tx : in std_logic_vector (1 downto 0);  
            data_tx_pl : out std_logic_vector (63 downto 0);  vc_write_tx_pl, 
            incr_tx_pl : out std_logic_vector (1 downto 0));
   end component;
   
   component output_register_vc_num2_vc_num_out2_3
      port( clk, rst : in std_logic;  data_tx : in std_logic_vector (63 downto 
            0);  vc_write_tx, incr_tx : in std_logic_vector (1 downto 0);  
            data_tx_pl : out std_logic_vector (63 downto 0);  vc_write_tx_pl, 
            incr_tx_pl : out std_logic_vector (1 downto 0));
   end component;
   
   component output_register_vc_num2_vc_num_out2_4
      port( clk, rst : in std_logic;  data_tx : in std_logic_vector (63 downto 
            0);  vc_write_tx, incr_tx : in std_logic_vector (1 downto 0);  
            data_tx_pl : out std_logic_vector (63 downto 0);  vc_write_tx_pl, 
            incr_tx_pl : out std_logic_vector (1 downto 0));
   end component;
   
   component output_register_vc_num2_vc_num_out2_5
      port( clk, rst : in std_logic;  data_tx : in std_logic_vector (63 downto 
            0);  vc_write_tx, incr_tx : in std_logic_vector (1 downto 0);  
            data_tx_pl : out std_logic_vector (63 downto 0);  vc_write_tx_pl, 
            incr_tx_pl : out std_logic_vector (1 downto 0));
   end component;
   
   component output_register_vc_num2_vc_num_out2_0
      port( clk, rst : in std_logic;  data_tx : in std_logic_vector (63 downto 
            0);  vc_write_tx, incr_tx : in std_logic_vector (1 downto 0);  
            data_tx_pl : out std_logic_vector (63 downto 0);  vc_write_tx_pl, 
            incr_tx_pl : out std_logic_vector (1 downto 0));
   end component;
   
   component output_register_vc_num1_vc_num_out1
      port( clk, rst : in std_logic;  data_tx : in std_logic_vector (63 downto 
            0);  vc_write_tx, incr_tx : in std_logic;  data_tx_pl : out 
            std_logic_vector (63 downto 0);  vc_write_tx_pl, incr_tx_pl : out 
            std_logic);
   end component;
   
   component crossbar_7_DXYU
      port( crossbar_in : in std_logic_vector (447 downto 0);  crossbar_ctrl : 
            in std_logic_vector (20 downto 0);  crossbar_out : out 
            std_logic_vector (447 downto 0));
   end component;
   
   component vc_input_buffer_2_0000000200000002_1
      port( clk, rst : in std_logic;  data_rx : in std_logic_vector (63 downto 
            0);  vc_write_rx, vc_transfer : in std_logic_vector (1 downto 0);  
            valid_data_vc : out std_logic_vector (1 downto 0);  data_transfer :
            out std_logic_vector (63 downto 0);  header : out std_logic_vector 
            (19 downto 0));
   end component;
   
   component vc_input_buffer_2_0000000200000002_2
      port( clk, rst : in std_logic;  data_rx : in std_logic_vector (63 downto 
            0);  vc_write_rx, vc_transfer : in std_logic_vector (1 downto 0);  
            valid_data_vc : out std_logic_vector (1 downto 0);  data_transfer :
            out std_logic_vector (63 downto 0);  header : out std_logic_vector 
            (19 downto 0));
   end component;
   
   component vc_input_buffer_2_0000000200000002_3
      port( clk, rst : in std_logic;  data_rx : in std_logic_vector (63 downto 
            0);  vc_write_rx, vc_transfer : in std_logic_vector (1 downto 0);  
            valid_data_vc : out std_logic_vector (1 downto 0);  data_transfer :
            out std_logic_vector (63 downto 0);  header : out std_logic_vector 
            (19 downto 0));
   end component;
   
   component vc_input_buffer_2_0000000200000002_4
      port( clk, rst : in std_logic;  data_rx : in std_logic_vector (63 downto 
            0);  vc_write_rx, vc_transfer : in std_logic_vector (1 downto 0);  
            valid_data_vc : out std_logic_vector (1 downto 0);  data_transfer :
            out std_logic_vector (63 downto 0);  header : out std_logic_vector 
            (19 downto 0));
   end component;
   
   component vc_input_buffer_2_0000000200000002_5
      port( clk, rst : in std_logic;  data_rx : in std_logic_vector (63 downto 
            0);  vc_write_rx, vc_transfer : in std_logic_vector (1 downto 0);  
            valid_data_vc : out std_logic_vector (1 downto 0);  data_transfer :
            out std_logic_vector (63 downto 0);  header : out std_logic_vector 
            (19 downto 0));
   end component;
   
   component vc_input_buffer_2_0000000200000002_0
      port( clk, rst : in std_logic;  data_rx : in std_logic_vector (63 downto 
            0);  vc_write_rx, vc_transfer : in std_logic_vector (1 downto 0);  
            valid_data_vc : out std_logic_vector (1 downto 0);  data_transfer :
            out std_logic_vector (63 downto 0);  header : out std_logic_vector 
            (19 downto 0));
   end component;
   
   component vc_input_buffer_1_0000000200000002
      port( clk, rst : in std_logic;  data_rx : in std_logic_vector (63 downto 
            0);  vc_write_rx, vc_transfer : in std_logic;  valid_data_vc : out 
            std_logic;  data_transfer : out std_logic_vector (63 downto 0);  
            header : out std_logic_vector (9 downto 0));
   end component;
   
   signal header_12_PACKET_LENGTH_3_port, header_12_PACKET_LENGTH_2_port, 
      header_12_PACKET_LENGTH_1_port, header_12_PACKET_LENGTH_0_port, 
      header_12_X_DEST_1_port, header_12_X_DEST_0_port, header_12_Y_DEST_1_port
      , header_12_Y_DEST_0_port, header_12_Z_DEST_1_port, 
      header_12_Z_DEST_0_port, header_11_PACKET_LENGTH_3_port, 
      header_11_PACKET_LENGTH_2_port, header_11_PACKET_LENGTH_1_port, 
      header_11_PACKET_LENGTH_0_port, header_11_X_DEST_1_port, 
      header_11_X_DEST_0_port, header_11_Y_DEST_1_port, header_11_Y_DEST_0_port
      , header_11_Z_DEST_1_port, header_11_Z_DEST_0_port, 
      header_10_PACKET_LENGTH_3_port, header_10_PACKET_LENGTH_2_port, 
      header_10_PACKET_LENGTH_1_port, header_10_PACKET_LENGTH_0_port, 
      header_10_X_DEST_1_port, header_10_X_DEST_0_port, header_10_Y_DEST_1_port
      , header_10_Y_DEST_0_port, header_10_Z_DEST_1_port, 
      header_10_Z_DEST_0_port, header_9_PACKET_LENGTH_3_port, 
      header_9_PACKET_LENGTH_2_port, header_9_PACKET_LENGTH_1_port, 
      header_9_PACKET_LENGTH_0_port, header_9_X_DEST_1_port, 
      header_9_X_DEST_0_port, header_9_Y_DEST_1_port, header_9_Y_DEST_0_port, 
      header_9_Z_DEST_1_port, header_9_Z_DEST_0_port, 
      header_8_PACKET_LENGTH_3_port, header_8_PACKET_LENGTH_2_port, 
      header_8_PACKET_LENGTH_1_port, header_8_PACKET_LENGTH_0_port, 
      header_8_X_DEST_1_port, header_8_X_DEST_0_port, header_8_Y_DEST_1_port, 
      header_8_Y_DEST_0_port, header_8_Z_DEST_1_port, header_8_Z_DEST_0_port, 
      header_7_PACKET_LENGTH_3_port, header_7_PACKET_LENGTH_2_port, 
      header_7_PACKET_LENGTH_1_port, header_7_PACKET_LENGTH_0_port, 
      header_7_X_DEST_1_port, header_7_X_DEST_0_port, header_7_Y_DEST_1_port, 
      header_7_Y_DEST_0_port, header_7_Z_DEST_1_port, header_7_Z_DEST_0_port, 
      header_6_PACKET_LENGTH_3_port, header_6_PACKET_LENGTH_2_port, 
      header_6_PACKET_LENGTH_1_port, header_6_PACKET_LENGTH_0_port, 
      header_6_X_DEST_1_port, header_6_X_DEST_0_port, header_6_Y_DEST_1_port, 
      header_6_Y_DEST_0_port, header_6_Z_DEST_1_port, header_6_Z_DEST_0_port, 
      header_5_PACKET_LENGTH_3_port, header_5_PACKET_LENGTH_2_port, 
      header_5_PACKET_LENGTH_1_port, header_5_PACKET_LENGTH_0_port, 
      header_5_X_DEST_1_port, header_5_X_DEST_0_port, header_5_Y_DEST_1_port, 
      header_5_Y_DEST_0_port, header_5_Z_DEST_1_port, header_5_Z_DEST_0_port, 
      header_4_PACKET_LENGTH_3_port, header_4_PACKET_LENGTH_2_port, 
      header_4_PACKET_LENGTH_1_port, header_4_PACKET_LENGTH_0_port, 
      header_4_X_DEST_1_port, header_4_X_DEST_0_port, header_4_Y_DEST_1_port, 
      header_4_Y_DEST_0_port, header_4_Z_DEST_1_port, header_4_Z_DEST_0_port, 
      header_3_PACKET_LENGTH_3_port, header_3_PACKET_LENGTH_2_port, 
      header_3_PACKET_LENGTH_1_port, header_3_PACKET_LENGTH_0_port, 
      header_3_X_DEST_1_port, header_3_X_DEST_0_port, header_3_Y_DEST_1_port, 
      header_3_Y_DEST_0_port, header_3_Z_DEST_1_port, header_3_Z_DEST_0_port, 
      header_2_PACKET_LENGTH_3_port, header_2_PACKET_LENGTH_2_port, 
      header_2_PACKET_LENGTH_1_port, header_2_PACKET_LENGTH_0_port, 
      header_2_X_DEST_1_port, header_2_X_DEST_0_port, header_2_Y_DEST_1_port, 
      header_2_Y_DEST_0_port, header_2_Z_DEST_1_port, header_2_Z_DEST_0_port, 
      header_1_PACKET_LENGTH_3_port, header_1_PACKET_LENGTH_2_port, 
      header_1_PACKET_LENGTH_1_port, header_1_PACKET_LENGTH_0_port, 
      header_1_X_DEST_1_port, header_1_X_DEST_0_port, header_1_Y_DEST_1_port, 
      header_1_Y_DEST_0_port, header_1_Z_DEST_1_port, header_1_Z_DEST_0_port, 
      header_0_PACKET_LENGTH_3_port, header_0_PACKET_LENGTH_2_port, 
      header_0_PACKET_LENGTH_1_port, header_0_PACKET_LENGTH_0_port, 
      header_0_X_DEST_1_port, header_0_X_DEST_0_port, header_0_Y_DEST_1_port, 
      header_0_Y_DEST_0_port, header_0_Z_DEST_1_port, header_0_Z_DEST_0_port, 
      data_transfer_6_63_port, data_transfer_6_62_port, data_transfer_6_61_port
      , data_transfer_6_60_port, data_transfer_6_59_port, 
      data_transfer_6_58_port, data_transfer_6_57_port, data_transfer_6_56_port
      , data_transfer_6_55_port, data_transfer_6_54_port, 
      data_transfer_6_53_port, data_transfer_6_52_port, data_transfer_6_51_port
      , data_transfer_6_50_port, data_transfer_6_49_port, 
      data_transfer_6_48_port, data_transfer_6_47_port, data_transfer_6_46_port
      , data_transfer_6_45_port, data_transfer_6_44_port, 
      data_transfer_6_43_port, data_transfer_6_42_port, data_transfer_6_41_port
      , data_transfer_6_40_port, data_transfer_6_39_port, 
      data_transfer_6_38_port, data_transfer_6_37_port, data_transfer_6_36_port
      , data_transfer_6_35_port, data_transfer_6_34_port, 
      data_transfer_6_33_port, data_transfer_6_32_port, data_transfer_6_31_port
      , data_transfer_6_30_port, data_transfer_6_29_port, 
      data_transfer_6_28_port, data_transfer_6_27_port, data_transfer_6_26_port
      , data_transfer_6_25_port, data_transfer_6_24_port, 
      data_transfer_6_23_port, data_transfer_6_22_port, data_transfer_6_21_port
      , data_transfer_6_20_port, data_transfer_6_19_port, 
      data_transfer_6_18_port, data_transfer_6_17_port, data_transfer_6_16_port
      , data_transfer_6_15_port, data_transfer_6_14_port, 
      data_transfer_6_13_port, data_transfer_6_12_port, data_transfer_6_11_port
      , data_transfer_6_10_port, data_transfer_6_9_port, data_transfer_6_8_port
      , data_transfer_6_7_port, data_transfer_6_6_port, data_transfer_6_5_port,
      data_transfer_6_4_port, data_transfer_6_3_port, data_transfer_6_2_port, 
      data_transfer_6_1_port, data_transfer_6_0_port, data_transfer_5_63_port, 
      data_transfer_5_62_port, data_transfer_5_61_port, data_transfer_5_60_port
      , data_transfer_5_59_port, data_transfer_5_58_port, 
      data_transfer_5_57_port, data_transfer_5_56_port, data_transfer_5_55_port
      , data_transfer_5_54_port, data_transfer_5_53_port, 
      data_transfer_5_52_port, data_transfer_5_51_port, data_transfer_5_50_port
      , data_transfer_5_49_port, data_transfer_5_48_port, 
      data_transfer_5_47_port, data_transfer_5_46_port, data_transfer_5_45_port
      , data_transfer_5_44_port, data_transfer_5_43_port, 
      data_transfer_5_42_port, data_transfer_5_41_port, data_transfer_5_40_port
      , data_transfer_5_39_port, data_transfer_5_38_port, 
      data_transfer_5_37_port, data_transfer_5_36_port, data_transfer_5_35_port
      , data_transfer_5_34_port, data_transfer_5_33_port, 
      data_transfer_5_32_port, data_transfer_5_31_port, data_transfer_5_30_port
      , data_transfer_5_29_port, data_transfer_5_28_port, 
      data_transfer_5_27_port, data_transfer_5_26_port, data_transfer_5_25_port
      , data_transfer_5_24_port, data_transfer_5_23_port, 
      data_transfer_5_22_port, data_transfer_5_21_port, data_transfer_5_20_port
      , data_transfer_5_19_port, data_transfer_5_18_port, 
      data_transfer_5_17_port, data_transfer_5_16_port, data_transfer_5_15_port
      , data_transfer_5_14_port, data_transfer_5_13_port, 
      data_transfer_5_12_port, data_transfer_5_11_port, data_transfer_5_10_port
      , data_transfer_5_9_port, data_transfer_5_8_port, data_transfer_5_7_port,
      data_transfer_5_6_port, data_transfer_5_5_port, data_transfer_5_4_port, 
      data_transfer_5_3_port, data_transfer_5_2_port, data_transfer_5_1_port, 
      data_transfer_5_0_port, data_transfer_4_63_port, data_transfer_4_62_port,
      data_transfer_4_61_port, data_transfer_4_60_port, data_transfer_4_59_port
      , data_transfer_4_58_port, data_transfer_4_57_port, 
      data_transfer_4_56_port, data_transfer_4_55_port, data_transfer_4_54_port
      , data_transfer_4_53_port, data_transfer_4_52_port, 
      data_transfer_4_51_port, data_transfer_4_50_port, data_transfer_4_49_port
      , data_transfer_4_48_port, data_transfer_4_47_port, 
      data_transfer_4_46_port, data_transfer_4_45_port, data_transfer_4_44_port
      , data_transfer_4_43_port, data_transfer_4_42_port, 
      data_transfer_4_41_port, data_transfer_4_40_port, data_transfer_4_39_port
      , data_transfer_4_38_port, data_transfer_4_37_port, 
      data_transfer_4_36_port, data_transfer_4_35_port, data_transfer_4_34_port
      , data_transfer_4_33_port, data_transfer_4_32_port, 
      data_transfer_4_31_port, data_transfer_4_30_port, data_transfer_4_29_port
      , data_transfer_4_28_port, data_transfer_4_27_port, 
      data_transfer_4_26_port, data_transfer_4_25_port, data_transfer_4_24_port
      , data_transfer_4_23_port, data_transfer_4_22_port, 
      data_transfer_4_21_port, data_transfer_4_20_port, data_transfer_4_19_port
      , data_transfer_4_18_port, data_transfer_4_17_port, 
      data_transfer_4_16_port, data_transfer_4_15_port, data_transfer_4_14_port
      , data_transfer_4_13_port, data_transfer_4_12_port, 
      data_transfer_4_11_port, data_transfer_4_10_port, data_transfer_4_9_port,
      data_transfer_4_8_port, data_transfer_4_7_port, data_transfer_4_6_port, 
      data_transfer_4_5_port, data_transfer_4_4_port, data_transfer_4_3_port, 
      data_transfer_4_2_port, data_transfer_4_1_port, data_transfer_4_0_port, 
      data_transfer_3_63_port, data_transfer_3_62_port, data_transfer_3_61_port
      , data_transfer_3_60_port, data_transfer_3_59_port, 
      data_transfer_3_58_port, data_transfer_3_57_port, data_transfer_3_56_port
      , data_transfer_3_55_port, data_transfer_3_54_port, 
      data_transfer_3_53_port, data_transfer_3_52_port, data_transfer_3_51_port
      , data_transfer_3_50_port, data_transfer_3_49_port, 
      data_transfer_3_48_port, data_transfer_3_47_port, data_transfer_3_46_port
      , data_transfer_3_45_port, data_transfer_3_44_port, 
      data_transfer_3_43_port, data_transfer_3_42_port, data_transfer_3_41_port
      , data_transfer_3_40_port, data_transfer_3_39_port, 
      data_transfer_3_38_port, data_transfer_3_37_port, data_transfer_3_36_port
      , data_transfer_3_35_port, data_transfer_3_34_port, 
      data_transfer_3_33_port, data_transfer_3_32_port, data_transfer_3_31_port
      , data_transfer_3_30_port, data_transfer_3_29_port, 
      data_transfer_3_28_port, data_transfer_3_27_port, data_transfer_3_26_port
      , data_transfer_3_25_port, data_transfer_3_24_port, 
      data_transfer_3_23_port, data_transfer_3_22_port, data_transfer_3_21_port
      , data_transfer_3_20_port, data_transfer_3_19_port, 
      data_transfer_3_18_port, data_transfer_3_17_port, data_transfer_3_16_port
      , data_transfer_3_15_port, data_transfer_3_14_port, 
      data_transfer_3_13_port, data_transfer_3_12_port, data_transfer_3_11_port
      , data_transfer_3_10_port, data_transfer_3_9_port, data_transfer_3_8_port
      , data_transfer_3_7_port, data_transfer_3_6_port, data_transfer_3_5_port,
      data_transfer_3_4_port, data_transfer_3_3_port, data_transfer_3_2_port, 
      data_transfer_3_1_port, data_transfer_3_0_port, data_transfer_2_63_port, 
      data_transfer_2_62_port, data_transfer_2_61_port, data_transfer_2_60_port
      , data_transfer_2_59_port, data_transfer_2_58_port, 
      data_transfer_2_57_port, data_transfer_2_56_port, data_transfer_2_55_port
      , data_transfer_2_54_port, data_transfer_2_53_port, 
      data_transfer_2_52_port, data_transfer_2_51_port, data_transfer_2_50_port
      , data_transfer_2_49_port, data_transfer_2_48_port, 
      data_transfer_2_47_port, data_transfer_2_46_port, data_transfer_2_45_port
      , data_transfer_2_44_port, data_transfer_2_43_port, 
      data_transfer_2_42_port, data_transfer_2_41_port, data_transfer_2_40_port
      , data_transfer_2_39_port, data_transfer_2_38_port, 
      data_transfer_2_37_port, data_transfer_2_36_port, data_transfer_2_35_port
      , data_transfer_2_34_port, data_transfer_2_33_port, 
      data_transfer_2_32_port, data_transfer_2_31_port, data_transfer_2_30_port
      , data_transfer_2_29_port, data_transfer_2_28_port, 
      data_transfer_2_27_port, data_transfer_2_26_port, data_transfer_2_25_port
      , data_transfer_2_24_port, data_transfer_2_23_port, 
      data_transfer_2_22_port, data_transfer_2_21_port, data_transfer_2_20_port
      , data_transfer_2_19_port, data_transfer_2_18_port, 
      data_transfer_2_17_port, data_transfer_2_16_port, data_transfer_2_15_port
      , data_transfer_2_14_port, data_transfer_2_13_port, 
      data_transfer_2_12_port, data_transfer_2_11_port, data_transfer_2_10_port
      , data_transfer_2_9_port, data_transfer_2_8_port, data_transfer_2_7_port,
      data_transfer_2_6_port, data_transfer_2_5_port, data_transfer_2_4_port, 
      data_transfer_2_3_port, data_transfer_2_2_port, data_transfer_2_1_port, 
      data_transfer_2_0_port, data_transfer_1_63_port, data_transfer_1_62_port,
      data_transfer_1_61_port, data_transfer_1_60_port, data_transfer_1_59_port
      , data_transfer_1_58_port, data_transfer_1_57_port, 
      data_transfer_1_56_port, data_transfer_1_55_port, data_transfer_1_54_port
      , data_transfer_1_53_port, data_transfer_1_52_port, 
      data_transfer_1_51_port, data_transfer_1_50_port, data_transfer_1_49_port
      , data_transfer_1_48_port, data_transfer_1_47_port, 
      data_transfer_1_46_port, data_transfer_1_45_port, data_transfer_1_44_port
      , data_transfer_1_43_port, data_transfer_1_42_port, 
      data_transfer_1_41_port, data_transfer_1_40_port, data_transfer_1_39_port
      , data_transfer_1_38_port, data_transfer_1_37_port, 
      data_transfer_1_36_port, data_transfer_1_35_port, data_transfer_1_34_port
      , data_transfer_1_33_port, data_transfer_1_32_port, 
      data_transfer_1_31_port, data_transfer_1_30_port, data_transfer_1_29_port
      , data_transfer_1_28_port, data_transfer_1_27_port, 
      data_transfer_1_26_port, data_transfer_1_25_port, data_transfer_1_24_port
      , data_transfer_1_23_port, data_transfer_1_22_port, 
      data_transfer_1_21_port, data_transfer_1_20_port, data_transfer_1_19_port
      , data_transfer_1_18_port, data_transfer_1_17_port, 
      data_transfer_1_16_port, data_transfer_1_15_port, data_transfer_1_14_port
      , data_transfer_1_13_port, data_transfer_1_12_port, 
      data_transfer_1_11_port, data_transfer_1_10_port, data_transfer_1_9_port,
      data_transfer_1_8_port, data_transfer_1_7_port, data_transfer_1_6_port, 
      data_transfer_1_5_port, data_transfer_1_4_port, data_transfer_1_3_port, 
      data_transfer_1_2_port, data_transfer_1_1_port, data_transfer_1_0_port, 
      data_transfer_0_63_port, data_transfer_0_62_port, data_transfer_0_61_port
      , data_transfer_0_60_port, data_transfer_0_59_port, 
      data_transfer_0_58_port, data_transfer_0_57_port, data_transfer_0_56_port
      , data_transfer_0_55_port, data_transfer_0_54_port, 
      data_transfer_0_53_port, data_transfer_0_52_port, data_transfer_0_51_port
      , data_transfer_0_50_port, data_transfer_0_49_port, 
      data_transfer_0_48_port, data_transfer_0_47_port, data_transfer_0_46_port
      , data_transfer_0_45_port, data_transfer_0_44_port, 
      data_transfer_0_43_port, data_transfer_0_42_port, data_transfer_0_41_port
      , data_transfer_0_40_port, data_transfer_0_39_port, 
      data_transfer_0_38_port, data_transfer_0_37_port, data_transfer_0_36_port
      , data_transfer_0_35_port, data_transfer_0_34_port, 
      data_transfer_0_33_port, data_transfer_0_32_port, data_transfer_0_31_port
      , data_transfer_0_30_port, data_transfer_0_29_port, 
      data_transfer_0_28_port, data_transfer_0_27_port, data_transfer_0_26_port
      , data_transfer_0_25_port, data_transfer_0_24_port, 
      data_transfer_0_23_port, data_transfer_0_22_port, data_transfer_0_21_port
      , data_transfer_0_20_port, data_transfer_0_19_port, 
      data_transfer_0_18_port, data_transfer_0_17_port, data_transfer_0_16_port
      , data_transfer_0_15_port, data_transfer_0_14_port, 
      data_transfer_0_13_port, data_transfer_0_12_port, data_transfer_0_11_port
      , data_transfer_0_10_port, data_transfer_0_9_port, data_transfer_0_8_port
      , data_transfer_0_7_port, data_transfer_0_6_port, data_transfer_0_5_port,
      data_transfer_0_4_port, data_transfer_0_3_port, data_transfer_0_2_port, 
      data_transfer_0_1_port, data_transfer_0_0_port, valid_data_vc_vec_12_port
      , valid_data_vc_vec_11_port, valid_data_vc_vec_10_port, 
      valid_data_vc_vec_9_port, valid_data_vc_vec_8_port, 
      valid_data_vc_vec_7_port, valid_data_vc_vec_6_port, 
      valid_data_vc_vec_5_port, valid_data_vc_vec_4_port, 
      valid_data_vc_vec_3_port, valid_data_vc_vec_2_port, 
      valid_data_vc_vec_1_port, valid_data_vc_vec_0_port, 
      vc_transfer_vec_12_port, vc_transfer_vec_11_port, vc_transfer_vec_10_port
      , vc_transfer_vec_9_port, vc_transfer_vec_8_port, vc_transfer_vec_7_port,
      vc_transfer_vec_6_port, vc_transfer_vec_5_port, vc_transfer_vec_4_port, 
      vc_transfer_vec_3_port, vc_transfer_vec_2_port, vc_transfer_vec_1_port, 
      vc_transfer_vec_0_port, crossbar_ctrl_20_port, crossbar_ctrl_19_port, 
      crossbar_ctrl_18_port, crossbar_ctrl_17_port, crossbar_ctrl_16_port, 
      crossbar_ctrl_15_port, crossbar_ctrl_14_port, crossbar_ctrl_13_port, 
      crossbar_ctrl_12_port, crossbar_ctrl_11_port, crossbar_ctrl_10_port, 
      crossbar_ctrl_9_port, crossbar_ctrl_8_port, crossbar_ctrl_7_port, 
      crossbar_ctrl_6_port, crossbar_ctrl_5_port, crossbar_ctrl_4_port, 
      crossbar_ctrl_3_port, crossbar_ctrl_2_port, crossbar_ctrl_1_port, 
      crossbar_ctrl_0_port, data_tx_6_63_port, data_tx_6_62_port, 
      data_tx_6_61_port, data_tx_6_60_port, data_tx_6_59_port, 
      data_tx_6_58_port, data_tx_6_57_port, data_tx_6_56_port, 
      data_tx_6_55_port, data_tx_6_54_port, data_tx_6_53_port, 
      data_tx_6_52_port, data_tx_6_51_port, data_tx_6_50_port, 
      data_tx_6_49_port, data_tx_6_48_port, data_tx_6_47_port, 
      data_tx_6_46_port, data_tx_6_45_port, data_tx_6_44_port, 
      data_tx_6_43_port, data_tx_6_42_port, data_tx_6_41_port, 
      data_tx_6_40_port, data_tx_6_39_port, data_tx_6_38_port, 
      data_tx_6_37_port, data_tx_6_36_port, data_tx_6_35_port, 
      data_tx_6_34_port, data_tx_6_33_port, data_tx_6_32_port, 
      data_tx_6_31_port, data_tx_6_30_port, data_tx_6_29_port, 
      data_tx_6_28_port, data_tx_6_27_port, data_tx_6_26_port, 
      data_tx_6_25_port, data_tx_6_24_port, data_tx_6_23_port, 
      data_tx_6_22_port, data_tx_6_21_port, data_tx_6_20_port, 
      data_tx_6_19_port, data_tx_6_18_port, data_tx_6_17_port, 
      data_tx_6_16_port, data_tx_6_15_port, data_tx_6_14_port, 
      data_tx_6_13_port, data_tx_6_12_port, data_tx_6_11_port, 
      data_tx_6_10_port, data_tx_6_9_port, data_tx_6_8_port, data_tx_6_7_port, 
      data_tx_6_6_port, data_tx_6_5_port, data_tx_6_4_port, data_tx_6_3_port, 
      data_tx_6_2_port, data_tx_6_1_port, data_tx_6_0_port, data_tx_5_63_port, 
      data_tx_5_62_port, data_tx_5_61_port, data_tx_5_60_port, 
      data_tx_5_59_port, data_tx_5_58_port, data_tx_5_57_port, 
      data_tx_5_56_port, data_tx_5_55_port, data_tx_5_54_port, 
      data_tx_5_53_port, data_tx_5_52_port, data_tx_5_51_port, 
      data_tx_5_50_port, data_tx_5_49_port, data_tx_5_48_port, 
      data_tx_5_47_port, data_tx_5_46_port, data_tx_5_45_port, 
      data_tx_5_44_port, data_tx_5_43_port, data_tx_5_42_port, 
      data_tx_5_41_port, data_tx_5_40_port, data_tx_5_39_port, 
      data_tx_5_38_port, data_tx_5_37_port, data_tx_5_36_port, 
      data_tx_5_35_port, data_tx_5_34_port, data_tx_5_33_port, 
      data_tx_5_32_port, data_tx_5_31_port, data_tx_5_30_port, 
      data_tx_5_29_port, data_tx_5_28_port, data_tx_5_27_port, 
      data_tx_5_26_port, data_tx_5_25_port, data_tx_5_24_port, 
      data_tx_5_23_port, data_tx_5_22_port, data_tx_5_21_port, 
      data_tx_5_20_port, data_tx_5_19_port, data_tx_5_18_port, 
      data_tx_5_17_port, data_tx_5_16_port, data_tx_5_15_port, 
      data_tx_5_14_port, data_tx_5_13_port, data_tx_5_12_port, 
      data_tx_5_11_port, data_tx_5_10_port, data_tx_5_9_port, data_tx_5_8_port,
      data_tx_5_7_port, data_tx_5_6_port, data_tx_5_5_port, data_tx_5_4_port, 
      data_tx_5_3_port, data_tx_5_2_port, data_tx_5_1_port, data_tx_5_0_port, 
      data_tx_4_63_port, data_tx_4_62_port, data_tx_4_61_port, 
      data_tx_4_60_port, data_tx_4_59_port, data_tx_4_58_port, 
      data_tx_4_57_port, data_tx_4_56_port, data_tx_4_55_port, 
      data_tx_4_54_port, data_tx_4_53_port, data_tx_4_52_port, 
      data_tx_4_51_port, data_tx_4_50_port, data_tx_4_49_port, 
      data_tx_4_48_port, data_tx_4_47_port, data_tx_4_46_port, 
      data_tx_4_45_port, data_tx_4_44_port, data_tx_4_43_port, 
      data_tx_4_42_port, data_tx_4_41_port, data_tx_4_40_port, 
      data_tx_4_39_port, data_tx_4_38_port, data_tx_4_37_port, 
      data_tx_4_36_port, data_tx_4_35_port, data_tx_4_34_port, 
      data_tx_4_33_port, data_tx_4_32_port, data_tx_4_31_port, 
      data_tx_4_30_port, data_tx_4_29_port, data_tx_4_28_port, 
      data_tx_4_27_port, data_tx_4_26_port, data_tx_4_25_port, 
      data_tx_4_24_port, data_tx_4_23_port, data_tx_4_22_port, 
      data_tx_4_21_port, data_tx_4_20_port, data_tx_4_19_port, 
      data_tx_4_18_port, data_tx_4_17_port, data_tx_4_16_port, 
      data_tx_4_15_port, data_tx_4_14_port, data_tx_4_13_port, 
      data_tx_4_12_port, data_tx_4_11_port, data_tx_4_10_port, data_tx_4_9_port
      , data_tx_4_8_port, data_tx_4_7_port, data_tx_4_6_port, data_tx_4_5_port,
      data_tx_4_4_port, data_tx_4_3_port, data_tx_4_2_port, data_tx_4_1_port, 
      data_tx_4_0_port, data_tx_3_63_port, data_tx_3_62_port, data_tx_3_61_port
      , data_tx_3_60_port, data_tx_3_59_port, data_tx_3_58_port, 
      data_tx_3_57_port, data_tx_3_56_port, data_tx_3_55_port, 
      data_tx_3_54_port, data_tx_3_53_port, data_tx_3_52_port, 
      data_tx_3_51_port, data_tx_3_50_port, data_tx_3_49_port, 
      data_tx_3_48_port, data_tx_3_47_port, data_tx_3_46_port, 
      data_tx_3_45_port, data_tx_3_44_port, data_tx_3_43_port, 
      data_tx_3_42_port, data_tx_3_41_port, data_tx_3_40_port, 
      data_tx_3_39_port, data_tx_3_38_port, data_tx_3_37_port, 
      data_tx_3_36_port, data_tx_3_35_port, data_tx_3_34_port, 
      data_tx_3_33_port, data_tx_3_32_port, data_tx_3_31_port, 
      data_tx_3_30_port, data_tx_3_29_port, data_tx_3_28_port, 
      data_tx_3_27_port, data_tx_3_26_port, data_tx_3_25_port, 
      data_tx_3_24_port, data_tx_3_23_port, data_tx_3_22_port, 
      data_tx_3_21_port, data_tx_3_20_port, data_tx_3_19_port, 
      data_tx_3_18_port, data_tx_3_17_port, data_tx_3_16_port, 
      data_tx_3_15_port, data_tx_3_14_port, data_tx_3_13_port, 
      data_tx_3_12_port, data_tx_3_11_port, data_tx_3_10_port, data_tx_3_9_port
      , data_tx_3_8_port, data_tx_3_7_port, data_tx_3_6_port, data_tx_3_5_port,
      data_tx_3_4_port, data_tx_3_3_port, data_tx_3_2_port, data_tx_3_1_port, 
      data_tx_3_0_port, data_tx_2_63_port, data_tx_2_62_port, data_tx_2_61_port
      , data_tx_2_60_port, data_tx_2_59_port, data_tx_2_58_port, 
      data_tx_2_57_port, data_tx_2_56_port, data_tx_2_55_port, 
      data_tx_2_54_port, data_tx_2_53_port, data_tx_2_52_port, 
      data_tx_2_51_port, data_tx_2_50_port, data_tx_2_49_port, 
      data_tx_2_48_port, data_tx_2_47_port, data_tx_2_46_port, 
      data_tx_2_45_port, data_tx_2_44_port, data_tx_2_43_port, 
      data_tx_2_42_port, data_tx_2_41_port, data_tx_2_40_port, 
      data_tx_2_39_port, data_tx_2_38_port, data_tx_2_37_port, 
      data_tx_2_36_port, data_tx_2_35_port, data_tx_2_34_port, 
      data_tx_2_33_port, data_tx_2_32_port, data_tx_2_31_port, 
      data_tx_2_30_port, data_tx_2_29_port, data_tx_2_28_port, 
      data_tx_2_27_port, data_tx_2_26_port, data_tx_2_25_port, 
      data_tx_2_24_port, data_tx_2_23_port, data_tx_2_22_port, 
      data_tx_2_21_port, data_tx_2_20_port, data_tx_2_19_port, 
      data_tx_2_18_port, data_tx_2_17_port, data_tx_2_16_port, 
      data_tx_2_15_port, data_tx_2_14_port, data_tx_2_13_port, 
      data_tx_2_12_port, data_tx_2_11_port, data_tx_2_10_port, data_tx_2_9_port
      , data_tx_2_8_port, data_tx_2_7_port, data_tx_2_6_port, data_tx_2_5_port,
      data_tx_2_4_port, data_tx_2_3_port, data_tx_2_2_port, data_tx_2_1_port, 
      data_tx_2_0_port, data_tx_1_63_port, data_tx_1_62_port, data_tx_1_61_port
      , data_tx_1_60_port, data_tx_1_59_port, data_tx_1_58_port, 
      data_tx_1_57_port, data_tx_1_56_port, data_tx_1_55_port, 
      data_tx_1_54_port, data_tx_1_53_port, data_tx_1_52_port, 
      data_tx_1_51_port, data_tx_1_50_port, data_tx_1_49_port, 
      data_tx_1_48_port, data_tx_1_47_port, data_tx_1_46_port, 
      data_tx_1_45_port, data_tx_1_44_port, data_tx_1_43_port, 
      data_tx_1_42_port, data_tx_1_41_port, data_tx_1_40_port, 
      data_tx_1_39_port, data_tx_1_38_port, data_tx_1_37_port, 
      data_tx_1_36_port, data_tx_1_35_port, data_tx_1_34_port, 
      data_tx_1_33_port, data_tx_1_32_port, data_tx_1_31_port, 
      data_tx_1_30_port, data_tx_1_29_port, data_tx_1_28_port, 
      data_tx_1_27_port, data_tx_1_26_port, data_tx_1_25_port, 
      data_tx_1_24_port, data_tx_1_23_port, data_tx_1_22_port, 
      data_tx_1_21_port, data_tx_1_20_port, data_tx_1_19_port, 
      data_tx_1_18_port, data_tx_1_17_port, data_tx_1_16_port, 
      data_tx_1_15_port, data_tx_1_14_port, data_tx_1_13_port, 
      data_tx_1_12_port, data_tx_1_11_port, data_tx_1_10_port, data_tx_1_9_port
      , data_tx_1_8_port, data_tx_1_7_port, data_tx_1_6_port, data_tx_1_5_port,
      data_tx_1_4_port, data_tx_1_3_port, data_tx_1_2_port, data_tx_1_1_port, 
      data_tx_1_0_port, data_tx_0_63_port, data_tx_0_62_port, data_tx_0_61_port
      , data_tx_0_60_port, data_tx_0_59_port, data_tx_0_58_port, 
      data_tx_0_57_port, data_tx_0_56_port, data_tx_0_55_port, 
      data_tx_0_54_port, data_tx_0_53_port, data_tx_0_52_port, 
      data_tx_0_51_port, data_tx_0_50_port, data_tx_0_49_port, 
      data_tx_0_48_port, data_tx_0_47_port, data_tx_0_46_port, 
      data_tx_0_45_port, data_tx_0_44_port, data_tx_0_43_port, 
      data_tx_0_42_port, data_tx_0_41_port, data_tx_0_40_port, 
      data_tx_0_39_port, data_tx_0_38_port, data_tx_0_37_port, 
      data_tx_0_36_port, data_tx_0_35_port, data_tx_0_34_port, 
      data_tx_0_33_port, data_tx_0_32_port, data_tx_0_31_port, 
      data_tx_0_30_port, data_tx_0_29_port, data_tx_0_28_port, 
      data_tx_0_27_port, data_tx_0_26_port, data_tx_0_25_port, 
      data_tx_0_24_port, data_tx_0_23_port, data_tx_0_22_port, 
      data_tx_0_21_port, data_tx_0_20_port, data_tx_0_19_port, 
      data_tx_0_18_port, data_tx_0_17_port, data_tx_0_16_port, 
      data_tx_0_15_port, data_tx_0_14_port, data_tx_0_13_port, 
      data_tx_0_12_port, data_tx_0_11_port, data_tx_0_10_port, data_tx_0_9_port
      , data_tx_0_8_port, data_tx_0_7_port, data_tx_0_6_port, data_tx_0_5_port,
      data_tx_0_4_port, data_tx_0_3_port, data_tx_0_2_port, data_tx_0_1_port, 
      data_tx_0_0_port, vc_write_tx_vec_12_port, vc_write_tx_vec_11_port, 
      vc_write_tx_vec_10_port, vc_write_tx_vec_9_port, vc_write_tx_vec_8_port, 
      vc_write_tx_vec_7_port, vc_write_tx_vec_6_port, vc_write_tx_vec_5_port, 
      vc_write_tx_vec_4_port, vc_write_tx_vec_3_port, vc_write_tx_vec_2_port, 
      vc_write_tx_vec_1_port, vc_write_tx_vec_0_port : std_logic;

begin
   
   vc_input_buffer_i_0 : vc_input_buffer_1_0000000200000002 port map( clk => 
                           clk, rst => rst, data_rx(63) => data_rx(0)(63), 
                           data_rx(62) => data_rx(0)(62), data_rx(61) => 
                           data_rx(0)(61), data_rx(60) => data_rx(0)(60), 
                           data_rx(59) => data_rx(0)(59), data_rx(58) => 
                           data_rx(0)(58), data_rx(57) => data_rx(0)(57), 
                           data_rx(56) => data_rx(0)(56), data_rx(55) => 
                           data_rx(0)(55), data_rx(54) => data_rx(0)(54), 
                           data_rx(53) => data_rx(0)(53), data_rx(52) => 
                           data_rx(0)(52), data_rx(51) => data_rx(0)(51), 
                           data_rx(50) => data_rx(0)(50), data_rx(49) => 
                           data_rx(0)(49), data_rx(48) => data_rx(0)(48), 
                           data_rx(47) => data_rx(0)(47), data_rx(46) => 
                           data_rx(0)(46), data_rx(45) => data_rx(0)(45), 
                           data_rx(44) => data_rx(0)(44), data_rx(43) => 
                           data_rx(0)(43), data_rx(42) => data_rx(0)(42), 
                           data_rx(41) => data_rx(0)(41), data_rx(40) => 
                           data_rx(0)(40), data_rx(39) => data_rx(0)(39), 
                           data_rx(38) => data_rx(0)(38), data_rx(37) => 
                           data_rx(0)(37), data_rx(36) => data_rx(0)(36), 
                           data_rx(35) => data_rx(0)(35), data_rx(34) => 
                           data_rx(0)(34), data_rx(33) => data_rx(0)(33), 
                           data_rx(32) => data_rx(0)(32), data_rx(31) => 
                           data_rx(0)(31), data_rx(30) => data_rx(0)(30), 
                           data_rx(29) => data_rx(0)(29), data_rx(28) => 
                           data_rx(0)(28), data_rx(27) => data_rx(0)(27), 
                           data_rx(26) => data_rx(0)(26), data_rx(25) => 
                           data_rx(0)(25), data_rx(24) => data_rx(0)(24), 
                           data_rx(23) => data_rx(0)(23), data_rx(22) => 
                           data_rx(0)(22), data_rx(21) => data_rx(0)(21), 
                           data_rx(20) => data_rx(0)(20), data_rx(19) => 
                           data_rx(0)(19), data_rx(18) => data_rx(0)(18), 
                           data_rx(17) => data_rx(0)(17), data_rx(16) => 
                           data_rx(0)(16), data_rx(15) => data_rx(0)(15), 
                           data_rx(14) => data_rx(0)(14), data_rx(13) => 
                           data_rx(0)(13), data_rx(12) => data_rx(0)(12), 
                           data_rx(11) => data_rx(0)(11), data_rx(10) => 
                           data_rx(0)(10), data_rx(9) => data_rx(0)(9), 
                           data_rx(8) => data_rx(0)(8), data_rx(7) => 
                           data_rx(0)(7), data_rx(6) => data_rx(0)(6), 
                           data_rx(5) => data_rx(0)(5), data_rx(4) => 
                           data_rx(0)(4), data_rx(3) => data_rx(0)(3), 
                           data_rx(2) => data_rx(0)(2), data_rx(1) => 
                           data_rx(0)(1), data_rx(0) => data_rx(0)(0), 
                           vc_write_rx => vc_write_rx_vec(0), vc_transfer => 
                           vc_transfer_vec_0_port, valid_data_vc => 
                           valid_data_vc_vec_0_port, data_transfer(63) => 
                           data_transfer_0_63_port, data_transfer(62) => 
                           data_transfer_0_62_port, data_transfer(61) => 
                           data_transfer_0_61_port, data_transfer(60) => 
                           data_transfer_0_60_port, data_transfer(59) => 
                           data_transfer_0_59_port, data_transfer(58) => 
                           data_transfer_0_58_port, data_transfer(57) => 
                           data_transfer_0_57_port, data_transfer(56) => 
                           data_transfer_0_56_port, data_transfer(55) => 
                           data_transfer_0_55_port, data_transfer(54) => 
                           data_transfer_0_54_port, data_transfer(53) => 
                           data_transfer_0_53_port, data_transfer(52) => 
                           data_transfer_0_52_port, data_transfer(51) => 
                           data_transfer_0_51_port, data_transfer(50) => 
                           data_transfer_0_50_port, data_transfer(49) => 
                           data_transfer_0_49_port, data_transfer(48) => 
                           data_transfer_0_48_port, data_transfer(47) => 
                           data_transfer_0_47_port, data_transfer(46) => 
                           data_transfer_0_46_port, data_transfer(45) => 
                           data_transfer_0_45_port, data_transfer(44) => 
                           data_transfer_0_44_port, data_transfer(43) => 
                           data_transfer_0_43_port, data_transfer(42) => 
                           data_transfer_0_42_port, data_transfer(41) => 
                           data_transfer_0_41_port, data_transfer(40) => 
                           data_transfer_0_40_port, data_transfer(39) => 
                           data_transfer_0_39_port, data_transfer(38) => 
                           data_transfer_0_38_port, data_transfer(37) => 
                           data_transfer_0_37_port, data_transfer(36) => 
                           data_transfer_0_36_port, data_transfer(35) => 
                           data_transfer_0_35_port, data_transfer(34) => 
                           data_transfer_0_34_port, data_transfer(33) => 
                           data_transfer_0_33_port, data_transfer(32) => 
                           data_transfer_0_32_port, data_transfer(31) => 
                           data_transfer_0_31_port, data_transfer(30) => 
                           data_transfer_0_30_port, data_transfer(29) => 
                           data_transfer_0_29_port, data_transfer(28) => 
                           data_transfer_0_28_port, data_transfer(27) => 
                           data_transfer_0_27_port, data_transfer(26) => 
                           data_transfer_0_26_port, data_transfer(25) => 
                           data_transfer_0_25_port, data_transfer(24) => 
                           data_transfer_0_24_port, data_transfer(23) => 
                           data_transfer_0_23_port, data_transfer(22) => 
                           data_transfer_0_22_port, data_transfer(21) => 
                           data_transfer_0_21_port, data_transfer(20) => 
                           data_transfer_0_20_port, data_transfer(19) => 
                           data_transfer_0_19_port, data_transfer(18) => 
                           data_transfer_0_18_port, data_transfer(17) => 
                           data_transfer_0_17_port, data_transfer(16) => 
                           data_transfer_0_16_port, data_transfer(15) => 
                           data_transfer_0_15_port, data_transfer(14) => 
                           data_transfer_0_14_port, data_transfer(13) => 
                           data_transfer_0_13_port, data_transfer(12) => 
                           data_transfer_0_12_port, data_transfer(11) => 
                           data_transfer_0_11_port, data_transfer(10) => 
                           data_transfer_0_10_port, data_transfer(9) => 
                           data_transfer_0_9_port, data_transfer(8) => 
                           data_transfer_0_8_port, data_transfer(7) => 
                           data_transfer_0_7_port, data_transfer(6) => 
                           data_transfer_0_6_port, data_transfer(5) => 
                           data_transfer_0_5_port, data_transfer(4) => 
                           data_transfer_0_4_port, data_transfer(3) => 
                           data_transfer_0_3_port, data_transfer(2) => 
                           data_transfer_0_2_port, data_transfer(1) => 
                           data_transfer_0_1_port, data_transfer(0) => 
                           data_transfer_0_0_port, header(9) => 
                           header_0_PACKET_LENGTH_3_port, header(8) => 
                           header_0_PACKET_LENGTH_2_port, header(7) => 
                           header_0_PACKET_LENGTH_1_port, header(6) => 
                           header_0_PACKET_LENGTH_0_port, header(5) => 
                           header_0_X_DEST_1_port, header(4) => 
                           header_0_X_DEST_0_port, header(3) => 
                           header_0_Y_DEST_1_port, header(2) => 
                           header_0_Y_DEST_0_port, header(1) => 
                           header_0_Z_DEST_1_port, header(0) => 
                           header_0_Z_DEST_0_port);
   vc_input_buffer_i_1 : vc_input_buffer_2_0000000200000002_0 port map( clk => 
                           clk, rst => rst, data_rx(63) => data_rx(1)(63), 
                           data_rx(62) => data_rx(1)(62), data_rx(61) => 
                           data_rx(1)(61), data_rx(60) => data_rx(1)(60), 
                           data_rx(59) => data_rx(1)(59), data_rx(58) => 
                           data_rx(1)(58), data_rx(57) => data_rx(1)(57), 
                           data_rx(56) => data_rx(1)(56), data_rx(55) => 
                           data_rx(1)(55), data_rx(54) => data_rx(1)(54), 
                           data_rx(53) => data_rx(1)(53), data_rx(52) => 
                           data_rx(1)(52), data_rx(51) => data_rx(1)(51), 
                           data_rx(50) => data_rx(1)(50), data_rx(49) => 
                           data_rx(1)(49), data_rx(48) => data_rx(1)(48), 
                           data_rx(47) => data_rx(1)(47), data_rx(46) => 
                           data_rx(1)(46), data_rx(45) => data_rx(1)(45), 
                           data_rx(44) => data_rx(1)(44), data_rx(43) => 
                           data_rx(1)(43), data_rx(42) => data_rx(1)(42), 
                           data_rx(41) => data_rx(1)(41), data_rx(40) => 
                           data_rx(1)(40), data_rx(39) => data_rx(1)(39), 
                           data_rx(38) => data_rx(1)(38), data_rx(37) => 
                           data_rx(1)(37), data_rx(36) => data_rx(1)(36), 
                           data_rx(35) => data_rx(1)(35), data_rx(34) => 
                           data_rx(1)(34), data_rx(33) => data_rx(1)(33), 
                           data_rx(32) => data_rx(1)(32), data_rx(31) => 
                           data_rx(1)(31), data_rx(30) => data_rx(1)(30), 
                           data_rx(29) => data_rx(1)(29), data_rx(28) => 
                           data_rx(1)(28), data_rx(27) => data_rx(1)(27), 
                           data_rx(26) => data_rx(1)(26), data_rx(25) => 
                           data_rx(1)(25), data_rx(24) => data_rx(1)(24), 
                           data_rx(23) => data_rx(1)(23), data_rx(22) => 
                           data_rx(1)(22), data_rx(21) => data_rx(1)(21), 
                           data_rx(20) => data_rx(1)(20), data_rx(19) => 
                           data_rx(1)(19), data_rx(18) => data_rx(1)(18), 
                           data_rx(17) => data_rx(1)(17), data_rx(16) => 
                           data_rx(1)(16), data_rx(15) => data_rx(1)(15), 
                           data_rx(14) => data_rx(1)(14), data_rx(13) => 
                           data_rx(1)(13), data_rx(12) => data_rx(1)(12), 
                           data_rx(11) => data_rx(1)(11), data_rx(10) => 
                           data_rx(1)(10), data_rx(9) => data_rx(1)(9), 
                           data_rx(8) => data_rx(1)(8), data_rx(7) => 
                           data_rx(1)(7), data_rx(6) => data_rx(1)(6), 
                           data_rx(5) => data_rx(1)(5), data_rx(4) => 
                           data_rx(1)(4), data_rx(3) => data_rx(1)(3), 
                           data_rx(2) => data_rx(1)(2), data_rx(1) => 
                           data_rx(1)(1), data_rx(0) => data_rx(1)(0), 
                           vc_write_rx(1) => vc_write_rx_vec(2), vc_write_rx(0)
                           => vc_write_rx_vec(1), vc_transfer(1) => 
                           vc_transfer_vec_2_port, vc_transfer(0) => 
                           vc_transfer_vec_1_port, valid_data_vc(1) => 
                           valid_data_vc_vec_2_port, valid_data_vc(0) => 
                           valid_data_vc_vec_1_port, data_transfer(63) => 
                           data_transfer_1_63_port, data_transfer(62) => 
                           data_transfer_1_62_port, data_transfer(61) => 
                           data_transfer_1_61_port, data_transfer(60) => 
                           data_transfer_1_60_port, data_transfer(59) => 
                           data_transfer_1_59_port, data_transfer(58) => 
                           data_transfer_1_58_port, data_transfer(57) => 
                           data_transfer_1_57_port, data_transfer(56) => 
                           data_transfer_1_56_port, data_transfer(55) => 
                           data_transfer_1_55_port, data_transfer(54) => 
                           data_transfer_1_54_port, data_transfer(53) => 
                           data_transfer_1_53_port, data_transfer(52) => 
                           data_transfer_1_52_port, data_transfer(51) => 
                           data_transfer_1_51_port, data_transfer(50) => 
                           data_transfer_1_50_port, data_transfer(49) => 
                           data_transfer_1_49_port, data_transfer(48) => 
                           data_transfer_1_48_port, data_transfer(47) => 
                           data_transfer_1_47_port, data_transfer(46) => 
                           data_transfer_1_46_port, data_transfer(45) => 
                           data_transfer_1_45_port, data_transfer(44) => 
                           data_transfer_1_44_port, data_transfer(43) => 
                           data_transfer_1_43_port, data_transfer(42) => 
                           data_transfer_1_42_port, data_transfer(41) => 
                           data_transfer_1_41_port, data_transfer(40) => 
                           data_transfer_1_40_port, data_transfer(39) => 
                           data_transfer_1_39_port, data_transfer(38) => 
                           data_transfer_1_38_port, data_transfer(37) => 
                           data_transfer_1_37_port, data_transfer(36) => 
                           data_transfer_1_36_port, data_transfer(35) => 
                           data_transfer_1_35_port, data_transfer(34) => 
                           data_transfer_1_34_port, data_transfer(33) => 
                           data_transfer_1_33_port, data_transfer(32) => 
                           data_transfer_1_32_port, data_transfer(31) => 
                           data_transfer_1_31_port, data_transfer(30) => 
                           data_transfer_1_30_port, data_transfer(29) => 
                           data_transfer_1_29_port, data_transfer(28) => 
                           data_transfer_1_28_port, data_transfer(27) => 
                           data_transfer_1_27_port, data_transfer(26) => 
                           data_transfer_1_26_port, data_transfer(25) => 
                           data_transfer_1_25_port, data_transfer(24) => 
                           data_transfer_1_24_port, data_transfer(23) => 
                           data_transfer_1_23_port, data_transfer(22) => 
                           data_transfer_1_22_port, data_transfer(21) => 
                           data_transfer_1_21_port, data_transfer(20) => 
                           data_transfer_1_20_port, data_transfer(19) => 
                           data_transfer_1_19_port, data_transfer(18) => 
                           data_transfer_1_18_port, data_transfer(17) => 
                           data_transfer_1_17_port, data_transfer(16) => 
                           data_transfer_1_16_port, data_transfer(15) => 
                           data_transfer_1_15_port, data_transfer(14) => 
                           data_transfer_1_14_port, data_transfer(13) => 
                           data_transfer_1_13_port, data_transfer(12) => 
                           data_transfer_1_12_port, data_transfer(11) => 
                           data_transfer_1_11_port, data_transfer(10) => 
                           data_transfer_1_10_port, data_transfer(9) => 
                           data_transfer_1_9_port, data_transfer(8) => 
                           data_transfer_1_8_port, data_transfer(7) => 
                           data_transfer_1_7_port, data_transfer(6) => 
                           data_transfer_1_6_port, data_transfer(5) => 
                           data_transfer_1_5_port, data_transfer(4) => 
                           data_transfer_1_4_port, data_transfer(3) => 
                           data_transfer_1_3_port, data_transfer(2) => 
                           data_transfer_1_2_port, data_transfer(1) => 
                           data_transfer_1_1_port, data_transfer(0) => 
                           data_transfer_1_0_port, header(19) => 
                           header_2_PACKET_LENGTH_3_port, header(18) => 
                           header_2_PACKET_LENGTH_2_port, header(17) => 
                           header_2_PACKET_LENGTH_1_port, header(16) => 
                           header_2_PACKET_LENGTH_0_port, header(15) => 
                           header_2_X_DEST_1_port, header(14) => 
                           header_2_X_DEST_0_port, header(13) => 
                           header_2_Y_DEST_1_port, header(12) => 
                           header_2_Y_DEST_0_port, header(11) => 
                           header_2_Z_DEST_1_port, header(10) => 
                           header_2_Z_DEST_0_port, header(9) => 
                           header_1_PACKET_LENGTH_3_port, header(8) => 
                           header_1_PACKET_LENGTH_2_port, header(7) => 
                           header_1_PACKET_LENGTH_1_port, header(6) => 
                           header_1_PACKET_LENGTH_0_port, header(5) => 
                           header_1_X_DEST_1_port, header(4) => 
                           header_1_X_DEST_0_port, header(3) => 
                           header_1_Y_DEST_1_port, header(2) => 
                           header_1_Y_DEST_0_port, header(1) => 
                           header_1_Z_DEST_1_port, header(0) => 
                           header_1_Z_DEST_0_port);
   vc_input_buffer_i_2 : vc_input_buffer_2_0000000200000002_5 port map( clk => 
                           clk, rst => rst, data_rx(63) => data_rx(2)(63), 
                           data_rx(62) => data_rx(2)(62), data_rx(61) => 
                           data_rx(2)(61), data_rx(60) => data_rx(2)(60), 
                           data_rx(59) => data_rx(2)(59), data_rx(58) => 
                           data_rx(2)(58), data_rx(57) => data_rx(2)(57), 
                           data_rx(56) => data_rx(2)(56), data_rx(55) => 
                           data_rx(2)(55), data_rx(54) => data_rx(2)(54), 
                           data_rx(53) => data_rx(2)(53), data_rx(52) => 
                           data_rx(2)(52), data_rx(51) => data_rx(2)(51), 
                           data_rx(50) => data_rx(2)(50), data_rx(49) => 
                           data_rx(2)(49), data_rx(48) => data_rx(2)(48), 
                           data_rx(47) => data_rx(2)(47), data_rx(46) => 
                           data_rx(2)(46), data_rx(45) => data_rx(2)(45), 
                           data_rx(44) => data_rx(2)(44), data_rx(43) => 
                           data_rx(2)(43), data_rx(42) => data_rx(2)(42), 
                           data_rx(41) => data_rx(2)(41), data_rx(40) => 
                           data_rx(2)(40), data_rx(39) => data_rx(2)(39), 
                           data_rx(38) => data_rx(2)(38), data_rx(37) => 
                           data_rx(2)(37), data_rx(36) => data_rx(2)(36), 
                           data_rx(35) => data_rx(2)(35), data_rx(34) => 
                           data_rx(2)(34), data_rx(33) => data_rx(2)(33), 
                           data_rx(32) => data_rx(2)(32), data_rx(31) => 
                           data_rx(2)(31), data_rx(30) => data_rx(2)(30), 
                           data_rx(29) => data_rx(2)(29), data_rx(28) => 
                           data_rx(2)(28), data_rx(27) => data_rx(2)(27), 
                           data_rx(26) => data_rx(2)(26), data_rx(25) => 
                           data_rx(2)(25), data_rx(24) => data_rx(2)(24), 
                           data_rx(23) => data_rx(2)(23), data_rx(22) => 
                           data_rx(2)(22), data_rx(21) => data_rx(2)(21), 
                           data_rx(20) => data_rx(2)(20), data_rx(19) => 
                           data_rx(2)(19), data_rx(18) => data_rx(2)(18), 
                           data_rx(17) => data_rx(2)(17), data_rx(16) => 
                           data_rx(2)(16), data_rx(15) => data_rx(2)(15), 
                           data_rx(14) => data_rx(2)(14), data_rx(13) => 
                           data_rx(2)(13), data_rx(12) => data_rx(2)(12), 
                           data_rx(11) => data_rx(2)(11), data_rx(10) => 
                           data_rx(2)(10), data_rx(9) => data_rx(2)(9), 
                           data_rx(8) => data_rx(2)(8), data_rx(7) => 
                           data_rx(2)(7), data_rx(6) => data_rx(2)(6), 
                           data_rx(5) => data_rx(2)(5), data_rx(4) => 
                           data_rx(2)(4), data_rx(3) => data_rx(2)(3), 
                           data_rx(2) => data_rx(2)(2), data_rx(1) => 
                           data_rx(2)(1), data_rx(0) => data_rx(2)(0), 
                           vc_write_rx(1) => vc_write_rx_vec(4), vc_write_rx(0)
                           => vc_write_rx_vec(3), vc_transfer(1) => 
                           vc_transfer_vec_4_port, vc_transfer(0) => 
                           vc_transfer_vec_3_port, valid_data_vc(1) => 
                           valid_data_vc_vec_4_port, valid_data_vc(0) => 
                           valid_data_vc_vec_3_port, data_transfer(63) => 
                           data_transfer_2_63_port, data_transfer(62) => 
                           data_transfer_2_62_port, data_transfer(61) => 
                           data_transfer_2_61_port, data_transfer(60) => 
                           data_transfer_2_60_port, data_transfer(59) => 
                           data_transfer_2_59_port, data_transfer(58) => 
                           data_transfer_2_58_port, data_transfer(57) => 
                           data_transfer_2_57_port, data_transfer(56) => 
                           data_transfer_2_56_port, data_transfer(55) => 
                           data_transfer_2_55_port, data_transfer(54) => 
                           data_transfer_2_54_port, data_transfer(53) => 
                           data_transfer_2_53_port, data_transfer(52) => 
                           data_transfer_2_52_port, data_transfer(51) => 
                           data_transfer_2_51_port, data_transfer(50) => 
                           data_transfer_2_50_port, data_transfer(49) => 
                           data_transfer_2_49_port, data_transfer(48) => 
                           data_transfer_2_48_port, data_transfer(47) => 
                           data_transfer_2_47_port, data_transfer(46) => 
                           data_transfer_2_46_port, data_transfer(45) => 
                           data_transfer_2_45_port, data_transfer(44) => 
                           data_transfer_2_44_port, data_transfer(43) => 
                           data_transfer_2_43_port, data_transfer(42) => 
                           data_transfer_2_42_port, data_transfer(41) => 
                           data_transfer_2_41_port, data_transfer(40) => 
                           data_transfer_2_40_port, data_transfer(39) => 
                           data_transfer_2_39_port, data_transfer(38) => 
                           data_transfer_2_38_port, data_transfer(37) => 
                           data_transfer_2_37_port, data_transfer(36) => 
                           data_transfer_2_36_port, data_transfer(35) => 
                           data_transfer_2_35_port, data_transfer(34) => 
                           data_transfer_2_34_port, data_transfer(33) => 
                           data_transfer_2_33_port, data_transfer(32) => 
                           data_transfer_2_32_port, data_transfer(31) => 
                           data_transfer_2_31_port, data_transfer(30) => 
                           data_transfer_2_30_port, data_transfer(29) => 
                           data_transfer_2_29_port, data_transfer(28) => 
                           data_transfer_2_28_port, data_transfer(27) => 
                           data_transfer_2_27_port, data_transfer(26) => 
                           data_transfer_2_26_port, data_transfer(25) => 
                           data_transfer_2_25_port, data_transfer(24) => 
                           data_transfer_2_24_port, data_transfer(23) => 
                           data_transfer_2_23_port, data_transfer(22) => 
                           data_transfer_2_22_port, data_transfer(21) => 
                           data_transfer_2_21_port, data_transfer(20) => 
                           data_transfer_2_20_port, data_transfer(19) => 
                           data_transfer_2_19_port, data_transfer(18) => 
                           data_transfer_2_18_port, data_transfer(17) => 
                           data_transfer_2_17_port, data_transfer(16) => 
                           data_transfer_2_16_port, data_transfer(15) => 
                           data_transfer_2_15_port, data_transfer(14) => 
                           data_transfer_2_14_port, data_transfer(13) => 
                           data_transfer_2_13_port, data_transfer(12) => 
                           data_transfer_2_12_port, data_transfer(11) => 
                           data_transfer_2_11_port, data_transfer(10) => 
                           data_transfer_2_10_port, data_transfer(9) => 
                           data_transfer_2_9_port, data_transfer(8) => 
                           data_transfer_2_8_port, data_transfer(7) => 
                           data_transfer_2_7_port, data_transfer(6) => 
                           data_transfer_2_6_port, data_transfer(5) => 
                           data_transfer_2_5_port, data_transfer(4) => 
                           data_transfer_2_4_port, data_transfer(3) => 
                           data_transfer_2_3_port, data_transfer(2) => 
                           data_transfer_2_2_port, data_transfer(1) => 
                           data_transfer_2_1_port, data_transfer(0) => 
                           data_transfer_2_0_port, header(19) => 
                           header_4_PACKET_LENGTH_3_port, header(18) => 
                           header_4_PACKET_LENGTH_2_port, header(17) => 
                           header_4_PACKET_LENGTH_1_port, header(16) => 
                           header_4_PACKET_LENGTH_0_port, header(15) => 
                           header_4_X_DEST_1_port, header(14) => 
                           header_4_X_DEST_0_port, header(13) => 
                           header_4_Y_DEST_1_port, header(12) => 
                           header_4_Y_DEST_0_port, header(11) => 
                           header_4_Z_DEST_1_port, header(10) => 
                           header_4_Z_DEST_0_port, header(9) => 
                           header_3_PACKET_LENGTH_3_port, header(8) => 
                           header_3_PACKET_LENGTH_2_port, header(7) => 
                           header_3_PACKET_LENGTH_1_port, header(6) => 
                           header_3_PACKET_LENGTH_0_port, header(5) => 
                           header_3_X_DEST_1_port, header(4) => 
                           header_3_X_DEST_0_port, header(3) => 
                           header_3_Y_DEST_1_port, header(2) => 
                           header_3_Y_DEST_0_port, header(1) => 
                           header_3_Z_DEST_1_port, header(0) => 
                           header_3_Z_DEST_0_port);
   vc_input_buffer_i_3 : vc_input_buffer_2_0000000200000002_4 port map( clk => 
                           clk, rst => rst, data_rx(63) => data_rx(3)(63), 
                           data_rx(62) => data_rx(3)(62), data_rx(61) => 
                           data_rx(3)(61), data_rx(60) => data_rx(3)(60), 
                           data_rx(59) => data_rx(3)(59), data_rx(58) => 
                           data_rx(3)(58), data_rx(57) => data_rx(3)(57), 
                           data_rx(56) => data_rx(3)(56), data_rx(55) => 
                           data_rx(3)(55), data_rx(54) => data_rx(3)(54), 
                           data_rx(53) => data_rx(3)(53), data_rx(52) => 
                           data_rx(3)(52), data_rx(51) => data_rx(3)(51), 
                           data_rx(50) => data_rx(3)(50), data_rx(49) => 
                           data_rx(3)(49), data_rx(48) => data_rx(3)(48), 
                           data_rx(47) => data_rx(3)(47), data_rx(46) => 
                           data_rx(3)(46), data_rx(45) => data_rx(3)(45), 
                           data_rx(44) => data_rx(3)(44), data_rx(43) => 
                           data_rx(3)(43), data_rx(42) => data_rx(3)(42), 
                           data_rx(41) => data_rx(3)(41), data_rx(40) => 
                           data_rx(3)(40), data_rx(39) => data_rx(3)(39), 
                           data_rx(38) => data_rx(3)(38), data_rx(37) => 
                           data_rx(3)(37), data_rx(36) => data_rx(3)(36), 
                           data_rx(35) => data_rx(3)(35), data_rx(34) => 
                           data_rx(3)(34), data_rx(33) => data_rx(3)(33), 
                           data_rx(32) => data_rx(3)(32), data_rx(31) => 
                           data_rx(3)(31), data_rx(30) => data_rx(3)(30), 
                           data_rx(29) => data_rx(3)(29), data_rx(28) => 
                           data_rx(3)(28), data_rx(27) => data_rx(3)(27), 
                           data_rx(26) => data_rx(3)(26), data_rx(25) => 
                           data_rx(3)(25), data_rx(24) => data_rx(3)(24), 
                           data_rx(23) => data_rx(3)(23), data_rx(22) => 
                           data_rx(3)(22), data_rx(21) => data_rx(3)(21), 
                           data_rx(20) => data_rx(3)(20), data_rx(19) => 
                           data_rx(3)(19), data_rx(18) => data_rx(3)(18), 
                           data_rx(17) => data_rx(3)(17), data_rx(16) => 
                           data_rx(3)(16), data_rx(15) => data_rx(3)(15), 
                           data_rx(14) => data_rx(3)(14), data_rx(13) => 
                           data_rx(3)(13), data_rx(12) => data_rx(3)(12), 
                           data_rx(11) => data_rx(3)(11), data_rx(10) => 
                           data_rx(3)(10), data_rx(9) => data_rx(3)(9), 
                           data_rx(8) => data_rx(3)(8), data_rx(7) => 
                           data_rx(3)(7), data_rx(6) => data_rx(3)(6), 
                           data_rx(5) => data_rx(3)(5), data_rx(4) => 
                           data_rx(3)(4), data_rx(3) => data_rx(3)(3), 
                           data_rx(2) => data_rx(3)(2), data_rx(1) => 
                           data_rx(3)(1), data_rx(0) => data_rx(3)(0), 
                           vc_write_rx(1) => vc_write_rx_vec(6), vc_write_rx(0)
                           => vc_write_rx_vec(5), vc_transfer(1) => 
                           vc_transfer_vec_6_port, vc_transfer(0) => 
                           vc_transfer_vec_5_port, valid_data_vc(1) => 
                           valid_data_vc_vec_6_port, valid_data_vc(0) => 
                           valid_data_vc_vec_5_port, data_transfer(63) => 
                           data_transfer_3_63_port, data_transfer(62) => 
                           data_transfer_3_62_port, data_transfer(61) => 
                           data_transfer_3_61_port, data_transfer(60) => 
                           data_transfer_3_60_port, data_transfer(59) => 
                           data_transfer_3_59_port, data_transfer(58) => 
                           data_transfer_3_58_port, data_transfer(57) => 
                           data_transfer_3_57_port, data_transfer(56) => 
                           data_transfer_3_56_port, data_transfer(55) => 
                           data_transfer_3_55_port, data_transfer(54) => 
                           data_transfer_3_54_port, data_transfer(53) => 
                           data_transfer_3_53_port, data_transfer(52) => 
                           data_transfer_3_52_port, data_transfer(51) => 
                           data_transfer_3_51_port, data_transfer(50) => 
                           data_transfer_3_50_port, data_transfer(49) => 
                           data_transfer_3_49_port, data_transfer(48) => 
                           data_transfer_3_48_port, data_transfer(47) => 
                           data_transfer_3_47_port, data_transfer(46) => 
                           data_transfer_3_46_port, data_transfer(45) => 
                           data_transfer_3_45_port, data_transfer(44) => 
                           data_transfer_3_44_port, data_transfer(43) => 
                           data_transfer_3_43_port, data_transfer(42) => 
                           data_transfer_3_42_port, data_transfer(41) => 
                           data_transfer_3_41_port, data_transfer(40) => 
                           data_transfer_3_40_port, data_transfer(39) => 
                           data_transfer_3_39_port, data_transfer(38) => 
                           data_transfer_3_38_port, data_transfer(37) => 
                           data_transfer_3_37_port, data_transfer(36) => 
                           data_transfer_3_36_port, data_transfer(35) => 
                           data_transfer_3_35_port, data_transfer(34) => 
                           data_transfer_3_34_port, data_transfer(33) => 
                           data_transfer_3_33_port, data_transfer(32) => 
                           data_transfer_3_32_port, data_transfer(31) => 
                           data_transfer_3_31_port, data_transfer(30) => 
                           data_transfer_3_30_port, data_transfer(29) => 
                           data_transfer_3_29_port, data_transfer(28) => 
                           data_transfer_3_28_port, data_transfer(27) => 
                           data_transfer_3_27_port, data_transfer(26) => 
                           data_transfer_3_26_port, data_transfer(25) => 
                           data_transfer_3_25_port, data_transfer(24) => 
                           data_transfer_3_24_port, data_transfer(23) => 
                           data_transfer_3_23_port, data_transfer(22) => 
                           data_transfer_3_22_port, data_transfer(21) => 
                           data_transfer_3_21_port, data_transfer(20) => 
                           data_transfer_3_20_port, data_transfer(19) => 
                           data_transfer_3_19_port, data_transfer(18) => 
                           data_transfer_3_18_port, data_transfer(17) => 
                           data_transfer_3_17_port, data_transfer(16) => 
                           data_transfer_3_16_port, data_transfer(15) => 
                           data_transfer_3_15_port, data_transfer(14) => 
                           data_transfer_3_14_port, data_transfer(13) => 
                           data_transfer_3_13_port, data_transfer(12) => 
                           data_transfer_3_12_port, data_transfer(11) => 
                           data_transfer_3_11_port, data_transfer(10) => 
                           data_transfer_3_10_port, data_transfer(9) => 
                           data_transfer_3_9_port, data_transfer(8) => 
                           data_transfer_3_8_port, data_transfer(7) => 
                           data_transfer_3_7_port, data_transfer(6) => 
                           data_transfer_3_6_port, data_transfer(5) => 
                           data_transfer_3_5_port, data_transfer(4) => 
                           data_transfer_3_4_port, data_transfer(3) => 
                           data_transfer_3_3_port, data_transfer(2) => 
                           data_transfer_3_2_port, data_transfer(1) => 
                           data_transfer_3_1_port, data_transfer(0) => 
                           data_transfer_3_0_port, header(19) => 
                           header_6_PACKET_LENGTH_3_port, header(18) => 
                           header_6_PACKET_LENGTH_2_port, header(17) => 
                           header_6_PACKET_LENGTH_1_port, header(16) => 
                           header_6_PACKET_LENGTH_0_port, header(15) => 
                           header_6_X_DEST_1_port, header(14) => 
                           header_6_X_DEST_0_port, header(13) => 
                           header_6_Y_DEST_1_port, header(12) => 
                           header_6_Y_DEST_0_port, header(11) => 
                           header_6_Z_DEST_1_port, header(10) => 
                           header_6_Z_DEST_0_port, header(9) => 
                           header_5_PACKET_LENGTH_3_port, header(8) => 
                           header_5_PACKET_LENGTH_2_port, header(7) => 
                           header_5_PACKET_LENGTH_1_port, header(6) => 
                           header_5_PACKET_LENGTH_0_port, header(5) => 
                           header_5_X_DEST_1_port, header(4) => 
                           header_5_X_DEST_0_port, header(3) => 
                           header_5_Y_DEST_1_port, header(2) => 
                           header_5_Y_DEST_0_port, header(1) => 
                           header_5_Z_DEST_1_port, header(0) => 
                           header_5_Z_DEST_0_port);
   vc_input_buffer_i_4 : vc_input_buffer_2_0000000200000002_3 port map( clk => 
                           clk, rst => rst, data_rx(63) => data_rx(4)(63), 
                           data_rx(62) => data_rx(4)(62), data_rx(61) => 
                           data_rx(4)(61), data_rx(60) => data_rx(4)(60), 
                           data_rx(59) => data_rx(4)(59), data_rx(58) => 
                           data_rx(4)(58), data_rx(57) => data_rx(4)(57), 
                           data_rx(56) => data_rx(4)(56), data_rx(55) => 
                           data_rx(4)(55), data_rx(54) => data_rx(4)(54), 
                           data_rx(53) => data_rx(4)(53), data_rx(52) => 
                           data_rx(4)(52), data_rx(51) => data_rx(4)(51), 
                           data_rx(50) => data_rx(4)(50), data_rx(49) => 
                           data_rx(4)(49), data_rx(48) => data_rx(4)(48), 
                           data_rx(47) => data_rx(4)(47), data_rx(46) => 
                           data_rx(4)(46), data_rx(45) => data_rx(4)(45), 
                           data_rx(44) => data_rx(4)(44), data_rx(43) => 
                           data_rx(4)(43), data_rx(42) => data_rx(4)(42), 
                           data_rx(41) => data_rx(4)(41), data_rx(40) => 
                           data_rx(4)(40), data_rx(39) => data_rx(4)(39), 
                           data_rx(38) => data_rx(4)(38), data_rx(37) => 
                           data_rx(4)(37), data_rx(36) => data_rx(4)(36), 
                           data_rx(35) => data_rx(4)(35), data_rx(34) => 
                           data_rx(4)(34), data_rx(33) => data_rx(4)(33), 
                           data_rx(32) => data_rx(4)(32), data_rx(31) => 
                           data_rx(4)(31), data_rx(30) => data_rx(4)(30), 
                           data_rx(29) => data_rx(4)(29), data_rx(28) => 
                           data_rx(4)(28), data_rx(27) => data_rx(4)(27), 
                           data_rx(26) => data_rx(4)(26), data_rx(25) => 
                           data_rx(4)(25), data_rx(24) => data_rx(4)(24), 
                           data_rx(23) => data_rx(4)(23), data_rx(22) => 
                           data_rx(4)(22), data_rx(21) => data_rx(4)(21), 
                           data_rx(20) => data_rx(4)(20), data_rx(19) => 
                           data_rx(4)(19), data_rx(18) => data_rx(4)(18), 
                           data_rx(17) => data_rx(4)(17), data_rx(16) => 
                           data_rx(4)(16), data_rx(15) => data_rx(4)(15), 
                           data_rx(14) => data_rx(4)(14), data_rx(13) => 
                           data_rx(4)(13), data_rx(12) => data_rx(4)(12), 
                           data_rx(11) => data_rx(4)(11), data_rx(10) => 
                           data_rx(4)(10), data_rx(9) => data_rx(4)(9), 
                           data_rx(8) => data_rx(4)(8), data_rx(7) => 
                           data_rx(4)(7), data_rx(6) => data_rx(4)(6), 
                           data_rx(5) => data_rx(4)(5), data_rx(4) => 
                           data_rx(4)(4), data_rx(3) => data_rx(4)(3), 
                           data_rx(2) => data_rx(4)(2), data_rx(1) => 
                           data_rx(4)(1), data_rx(0) => data_rx(4)(0), 
                           vc_write_rx(1) => vc_write_rx_vec(8), vc_write_rx(0)
                           => vc_write_rx_vec(7), vc_transfer(1) => 
                           vc_transfer_vec_8_port, vc_transfer(0) => 
                           vc_transfer_vec_7_port, valid_data_vc(1) => 
                           valid_data_vc_vec_8_port, valid_data_vc(0) => 
                           valid_data_vc_vec_7_port, data_transfer(63) => 
                           data_transfer_4_63_port, data_transfer(62) => 
                           data_transfer_4_62_port, data_transfer(61) => 
                           data_transfer_4_61_port, data_transfer(60) => 
                           data_transfer_4_60_port, data_transfer(59) => 
                           data_transfer_4_59_port, data_transfer(58) => 
                           data_transfer_4_58_port, data_transfer(57) => 
                           data_transfer_4_57_port, data_transfer(56) => 
                           data_transfer_4_56_port, data_transfer(55) => 
                           data_transfer_4_55_port, data_transfer(54) => 
                           data_transfer_4_54_port, data_transfer(53) => 
                           data_transfer_4_53_port, data_transfer(52) => 
                           data_transfer_4_52_port, data_transfer(51) => 
                           data_transfer_4_51_port, data_transfer(50) => 
                           data_transfer_4_50_port, data_transfer(49) => 
                           data_transfer_4_49_port, data_transfer(48) => 
                           data_transfer_4_48_port, data_transfer(47) => 
                           data_transfer_4_47_port, data_transfer(46) => 
                           data_transfer_4_46_port, data_transfer(45) => 
                           data_transfer_4_45_port, data_transfer(44) => 
                           data_transfer_4_44_port, data_transfer(43) => 
                           data_transfer_4_43_port, data_transfer(42) => 
                           data_transfer_4_42_port, data_transfer(41) => 
                           data_transfer_4_41_port, data_transfer(40) => 
                           data_transfer_4_40_port, data_transfer(39) => 
                           data_transfer_4_39_port, data_transfer(38) => 
                           data_transfer_4_38_port, data_transfer(37) => 
                           data_transfer_4_37_port, data_transfer(36) => 
                           data_transfer_4_36_port, data_transfer(35) => 
                           data_transfer_4_35_port, data_transfer(34) => 
                           data_transfer_4_34_port, data_transfer(33) => 
                           data_transfer_4_33_port, data_transfer(32) => 
                           data_transfer_4_32_port, data_transfer(31) => 
                           data_transfer_4_31_port, data_transfer(30) => 
                           data_transfer_4_30_port, data_transfer(29) => 
                           data_transfer_4_29_port, data_transfer(28) => 
                           data_transfer_4_28_port, data_transfer(27) => 
                           data_transfer_4_27_port, data_transfer(26) => 
                           data_transfer_4_26_port, data_transfer(25) => 
                           data_transfer_4_25_port, data_transfer(24) => 
                           data_transfer_4_24_port, data_transfer(23) => 
                           data_transfer_4_23_port, data_transfer(22) => 
                           data_transfer_4_22_port, data_transfer(21) => 
                           data_transfer_4_21_port, data_transfer(20) => 
                           data_transfer_4_20_port, data_transfer(19) => 
                           data_transfer_4_19_port, data_transfer(18) => 
                           data_transfer_4_18_port, data_transfer(17) => 
                           data_transfer_4_17_port, data_transfer(16) => 
                           data_transfer_4_16_port, data_transfer(15) => 
                           data_transfer_4_15_port, data_transfer(14) => 
                           data_transfer_4_14_port, data_transfer(13) => 
                           data_transfer_4_13_port, data_transfer(12) => 
                           data_transfer_4_12_port, data_transfer(11) => 
                           data_transfer_4_11_port, data_transfer(10) => 
                           data_transfer_4_10_port, data_transfer(9) => 
                           data_transfer_4_9_port, data_transfer(8) => 
                           data_transfer_4_8_port, data_transfer(7) => 
                           data_transfer_4_7_port, data_transfer(6) => 
                           data_transfer_4_6_port, data_transfer(5) => 
                           data_transfer_4_5_port, data_transfer(4) => 
                           data_transfer_4_4_port, data_transfer(3) => 
                           data_transfer_4_3_port, data_transfer(2) => 
                           data_transfer_4_2_port, data_transfer(1) => 
                           data_transfer_4_1_port, data_transfer(0) => 
                           data_transfer_4_0_port, header(19) => 
                           header_8_PACKET_LENGTH_3_port, header(18) => 
                           header_8_PACKET_LENGTH_2_port, header(17) => 
                           header_8_PACKET_LENGTH_1_port, header(16) => 
                           header_8_PACKET_LENGTH_0_port, header(15) => 
                           header_8_X_DEST_1_port, header(14) => 
                           header_8_X_DEST_0_port, header(13) => 
                           header_8_Y_DEST_1_port, header(12) => 
                           header_8_Y_DEST_0_port, header(11) => 
                           header_8_Z_DEST_1_port, header(10) => 
                           header_8_Z_DEST_0_port, header(9) => 
                           header_7_PACKET_LENGTH_3_port, header(8) => 
                           header_7_PACKET_LENGTH_2_port, header(7) => 
                           header_7_PACKET_LENGTH_1_port, header(6) => 
                           header_7_PACKET_LENGTH_0_port, header(5) => 
                           header_7_X_DEST_1_port, header(4) => 
                           header_7_X_DEST_0_port, header(3) => 
                           header_7_Y_DEST_1_port, header(2) => 
                           header_7_Y_DEST_0_port, header(1) => 
                           header_7_Z_DEST_1_port, header(0) => 
                           header_7_Z_DEST_0_port);
   vc_input_buffer_i_5 : vc_input_buffer_2_0000000200000002_2 port map( clk => 
                           clk, rst => rst, data_rx(63) => data_rx(5)(63), 
                           data_rx(62) => data_rx(5)(62), data_rx(61) => 
                           data_rx(5)(61), data_rx(60) => data_rx(5)(60), 
                           data_rx(59) => data_rx(5)(59), data_rx(58) => 
                           data_rx(5)(58), data_rx(57) => data_rx(5)(57), 
                           data_rx(56) => data_rx(5)(56), data_rx(55) => 
                           data_rx(5)(55), data_rx(54) => data_rx(5)(54), 
                           data_rx(53) => data_rx(5)(53), data_rx(52) => 
                           data_rx(5)(52), data_rx(51) => data_rx(5)(51), 
                           data_rx(50) => data_rx(5)(50), data_rx(49) => 
                           data_rx(5)(49), data_rx(48) => data_rx(5)(48), 
                           data_rx(47) => data_rx(5)(47), data_rx(46) => 
                           data_rx(5)(46), data_rx(45) => data_rx(5)(45), 
                           data_rx(44) => data_rx(5)(44), data_rx(43) => 
                           data_rx(5)(43), data_rx(42) => data_rx(5)(42), 
                           data_rx(41) => data_rx(5)(41), data_rx(40) => 
                           data_rx(5)(40), data_rx(39) => data_rx(5)(39), 
                           data_rx(38) => data_rx(5)(38), data_rx(37) => 
                           data_rx(5)(37), data_rx(36) => data_rx(5)(36), 
                           data_rx(35) => data_rx(5)(35), data_rx(34) => 
                           data_rx(5)(34), data_rx(33) => data_rx(5)(33), 
                           data_rx(32) => data_rx(5)(32), data_rx(31) => 
                           data_rx(5)(31), data_rx(30) => data_rx(5)(30), 
                           data_rx(29) => data_rx(5)(29), data_rx(28) => 
                           data_rx(5)(28), data_rx(27) => data_rx(5)(27), 
                           data_rx(26) => data_rx(5)(26), data_rx(25) => 
                           data_rx(5)(25), data_rx(24) => data_rx(5)(24), 
                           data_rx(23) => data_rx(5)(23), data_rx(22) => 
                           data_rx(5)(22), data_rx(21) => data_rx(5)(21), 
                           data_rx(20) => data_rx(5)(20), data_rx(19) => 
                           data_rx(5)(19), data_rx(18) => data_rx(5)(18), 
                           data_rx(17) => data_rx(5)(17), data_rx(16) => 
                           data_rx(5)(16), data_rx(15) => data_rx(5)(15), 
                           data_rx(14) => data_rx(5)(14), data_rx(13) => 
                           data_rx(5)(13), data_rx(12) => data_rx(5)(12), 
                           data_rx(11) => data_rx(5)(11), data_rx(10) => 
                           data_rx(5)(10), data_rx(9) => data_rx(5)(9), 
                           data_rx(8) => data_rx(5)(8), data_rx(7) => 
                           data_rx(5)(7), data_rx(6) => data_rx(5)(6), 
                           data_rx(5) => data_rx(5)(5), data_rx(4) => 
                           data_rx(5)(4), data_rx(3) => data_rx(5)(3), 
                           data_rx(2) => data_rx(5)(2), data_rx(1) => 
                           data_rx(5)(1), data_rx(0) => data_rx(5)(0), 
                           vc_write_rx(1) => vc_write_rx_vec(10), 
                           vc_write_rx(0) => vc_write_rx_vec(9), vc_transfer(1)
                           => vc_transfer_vec_10_port, vc_transfer(0) => 
                           vc_transfer_vec_9_port, valid_data_vc(1) => 
                           valid_data_vc_vec_10_port, valid_data_vc(0) => 
                           valid_data_vc_vec_9_port, data_transfer(63) => 
                           data_transfer_5_63_port, data_transfer(62) => 
                           data_transfer_5_62_port, data_transfer(61) => 
                           data_transfer_5_61_port, data_transfer(60) => 
                           data_transfer_5_60_port, data_transfer(59) => 
                           data_transfer_5_59_port, data_transfer(58) => 
                           data_transfer_5_58_port, data_transfer(57) => 
                           data_transfer_5_57_port, data_transfer(56) => 
                           data_transfer_5_56_port, data_transfer(55) => 
                           data_transfer_5_55_port, data_transfer(54) => 
                           data_transfer_5_54_port, data_transfer(53) => 
                           data_transfer_5_53_port, data_transfer(52) => 
                           data_transfer_5_52_port, data_transfer(51) => 
                           data_transfer_5_51_port, data_transfer(50) => 
                           data_transfer_5_50_port, data_transfer(49) => 
                           data_transfer_5_49_port, data_transfer(48) => 
                           data_transfer_5_48_port, data_transfer(47) => 
                           data_transfer_5_47_port, data_transfer(46) => 
                           data_transfer_5_46_port, data_transfer(45) => 
                           data_transfer_5_45_port, data_transfer(44) => 
                           data_transfer_5_44_port, data_transfer(43) => 
                           data_transfer_5_43_port, data_transfer(42) => 
                           data_transfer_5_42_port, data_transfer(41) => 
                           data_transfer_5_41_port, data_transfer(40) => 
                           data_transfer_5_40_port, data_transfer(39) => 
                           data_transfer_5_39_port, data_transfer(38) => 
                           data_transfer_5_38_port, data_transfer(37) => 
                           data_transfer_5_37_port, data_transfer(36) => 
                           data_transfer_5_36_port, data_transfer(35) => 
                           data_transfer_5_35_port, data_transfer(34) => 
                           data_transfer_5_34_port, data_transfer(33) => 
                           data_transfer_5_33_port, data_transfer(32) => 
                           data_transfer_5_32_port, data_transfer(31) => 
                           data_transfer_5_31_port, data_transfer(30) => 
                           data_transfer_5_30_port, data_transfer(29) => 
                           data_transfer_5_29_port, data_transfer(28) => 
                           data_transfer_5_28_port, data_transfer(27) => 
                           data_transfer_5_27_port, data_transfer(26) => 
                           data_transfer_5_26_port, data_transfer(25) => 
                           data_transfer_5_25_port, data_transfer(24) => 
                           data_transfer_5_24_port, data_transfer(23) => 
                           data_transfer_5_23_port, data_transfer(22) => 
                           data_transfer_5_22_port, data_transfer(21) => 
                           data_transfer_5_21_port, data_transfer(20) => 
                           data_transfer_5_20_port, data_transfer(19) => 
                           data_transfer_5_19_port, data_transfer(18) => 
                           data_transfer_5_18_port, data_transfer(17) => 
                           data_transfer_5_17_port, data_transfer(16) => 
                           data_transfer_5_16_port, data_transfer(15) => 
                           data_transfer_5_15_port, data_transfer(14) => 
                           data_transfer_5_14_port, data_transfer(13) => 
                           data_transfer_5_13_port, data_transfer(12) => 
                           data_transfer_5_12_port, data_transfer(11) => 
                           data_transfer_5_11_port, data_transfer(10) => 
                           data_transfer_5_10_port, data_transfer(9) => 
                           data_transfer_5_9_port, data_transfer(8) => 
                           data_transfer_5_8_port, data_transfer(7) => 
                           data_transfer_5_7_port, data_transfer(6) => 
                           data_transfer_5_6_port, data_transfer(5) => 
                           data_transfer_5_5_port, data_transfer(4) => 
                           data_transfer_5_4_port, data_transfer(3) => 
                           data_transfer_5_3_port, data_transfer(2) => 
                           data_transfer_5_2_port, data_transfer(1) => 
                           data_transfer_5_1_port, data_transfer(0) => 
                           data_transfer_5_0_port, header(19) => 
                           header_10_PACKET_LENGTH_3_port, header(18) => 
                           header_10_PACKET_LENGTH_2_port, header(17) => 
                           header_10_PACKET_LENGTH_1_port, header(16) => 
                           header_10_PACKET_LENGTH_0_port, header(15) => 
                           header_10_X_DEST_1_port, header(14) => 
                           header_10_X_DEST_0_port, header(13) => 
                           header_10_Y_DEST_1_port, header(12) => 
                           header_10_Y_DEST_0_port, header(11) => 
                           header_10_Z_DEST_1_port, header(10) => 
                           header_10_Z_DEST_0_port, header(9) => 
                           header_9_PACKET_LENGTH_3_port, header(8) => 
                           header_9_PACKET_LENGTH_2_port, header(7) => 
                           header_9_PACKET_LENGTH_1_port, header(6) => 
                           header_9_PACKET_LENGTH_0_port, header(5) => 
                           header_9_X_DEST_1_port, header(4) => 
                           header_9_X_DEST_0_port, header(3) => 
                           header_9_Y_DEST_1_port, header(2) => 
                           header_9_Y_DEST_0_port, header(1) => 
                           header_9_Z_DEST_1_port, header(0) => 
                           header_9_Z_DEST_0_port);
   vc_input_buffer_i_6 : vc_input_buffer_2_0000000200000002_1 port map( clk => 
                           clk, rst => rst, data_rx(63) => data_rx(6)(63), 
                           data_rx(62) => data_rx(6)(62), data_rx(61) => 
                           data_rx(6)(61), data_rx(60) => data_rx(6)(60), 
                           data_rx(59) => data_rx(6)(59), data_rx(58) => 
                           data_rx(6)(58), data_rx(57) => data_rx(6)(57), 
                           data_rx(56) => data_rx(6)(56), data_rx(55) => 
                           data_rx(6)(55), data_rx(54) => data_rx(6)(54), 
                           data_rx(53) => data_rx(6)(53), data_rx(52) => 
                           data_rx(6)(52), data_rx(51) => data_rx(6)(51), 
                           data_rx(50) => data_rx(6)(50), data_rx(49) => 
                           data_rx(6)(49), data_rx(48) => data_rx(6)(48), 
                           data_rx(47) => data_rx(6)(47), data_rx(46) => 
                           data_rx(6)(46), data_rx(45) => data_rx(6)(45), 
                           data_rx(44) => data_rx(6)(44), data_rx(43) => 
                           data_rx(6)(43), data_rx(42) => data_rx(6)(42), 
                           data_rx(41) => data_rx(6)(41), data_rx(40) => 
                           data_rx(6)(40), data_rx(39) => data_rx(6)(39), 
                           data_rx(38) => data_rx(6)(38), data_rx(37) => 
                           data_rx(6)(37), data_rx(36) => data_rx(6)(36), 
                           data_rx(35) => data_rx(6)(35), data_rx(34) => 
                           data_rx(6)(34), data_rx(33) => data_rx(6)(33), 
                           data_rx(32) => data_rx(6)(32), data_rx(31) => 
                           data_rx(6)(31), data_rx(30) => data_rx(6)(30), 
                           data_rx(29) => data_rx(6)(29), data_rx(28) => 
                           data_rx(6)(28), data_rx(27) => data_rx(6)(27), 
                           data_rx(26) => data_rx(6)(26), data_rx(25) => 
                           data_rx(6)(25), data_rx(24) => data_rx(6)(24), 
                           data_rx(23) => data_rx(6)(23), data_rx(22) => 
                           data_rx(6)(22), data_rx(21) => data_rx(6)(21), 
                           data_rx(20) => data_rx(6)(20), data_rx(19) => 
                           data_rx(6)(19), data_rx(18) => data_rx(6)(18), 
                           data_rx(17) => data_rx(6)(17), data_rx(16) => 
                           data_rx(6)(16), data_rx(15) => data_rx(6)(15), 
                           data_rx(14) => data_rx(6)(14), data_rx(13) => 
                           data_rx(6)(13), data_rx(12) => data_rx(6)(12), 
                           data_rx(11) => data_rx(6)(11), data_rx(10) => 
                           data_rx(6)(10), data_rx(9) => data_rx(6)(9), 
                           data_rx(8) => data_rx(6)(8), data_rx(7) => 
                           data_rx(6)(7), data_rx(6) => data_rx(6)(6), 
                           data_rx(5) => data_rx(6)(5), data_rx(4) => 
                           data_rx(6)(4), data_rx(3) => data_rx(6)(3), 
                           data_rx(2) => data_rx(6)(2), data_rx(1) => 
                           data_rx(6)(1), data_rx(0) => data_rx(6)(0), 
                           vc_write_rx(1) => vc_write_rx_vec(12), 
                           vc_write_rx(0) => vc_write_rx_vec(11), 
                           vc_transfer(1) => vc_transfer_vec_12_port, 
                           vc_transfer(0) => vc_transfer_vec_11_port, 
                           valid_data_vc(1) => valid_data_vc_vec_12_port, 
                           valid_data_vc(0) => valid_data_vc_vec_11_port, 
                           data_transfer(63) => data_transfer_6_63_port, 
                           data_transfer(62) => data_transfer_6_62_port, 
                           data_transfer(61) => data_transfer_6_61_port, 
                           data_transfer(60) => data_transfer_6_60_port, 
                           data_transfer(59) => data_transfer_6_59_port, 
                           data_transfer(58) => data_transfer_6_58_port, 
                           data_transfer(57) => data_transfer_6_57_port, 
                           data_transfer(56) => data_transfer_6_56_port, 
                           data_transfer(55) => data_transfer_6_55_port, 
                           data_transfer(54) => data_transfer_6_54_port, 
                           data_transfer(53) => data_transfer_6_53_port, 
                           data_transfer(52) => data_transfer_6_52_port, 
                           data_transfer(51) => data_transfer_6_51_port, 
                           data_transfer(50) => data_transfer_6_50_port, 
                           data_transfer(49) => data_transfer_6_49_port, 
                           data_transfer(48) => data_transfer_6_48_port, 
                           data_transfer(47) => data_transfer_6_47_port, 
                           data_transfer(46) => data_transfer_6_46_port, 
                           data_transfer(45) => data_transfer_6_45_port, 
                           data_transfer(44) => data_transfer_6_44_port, 
                           data_transfer(43) => data_transfer_6_43_port, 
                           data_transfer(42) => data_transfer_6_42_port, 
                           data_transfer(41) => data_transfer_6_41_port, 
                           data_transfer(40) => data_transfer_6_40_port, 
                           data_transfer(39) => data_transfer_6_39_port, 
                           data_transfer(38) => data_transfer_6_38_port, 
                           data_transfer(37) => data_transfer_6_37_port, 
                           data_transfer(36) => data_transfer_6_36_port, 
                           data_transfer(35) => data_transfer_6_35_port, 
                           data_transfer(34) => data_transfer_6_34_port, 
                           data_transfer(33) => data_transfer_6_33_port, 
                           data_transfer(32) => data_transfer_6_32_port, 
                           data_transfer(31) => data_transfer_6_31_port, 
                           data_transfer(30) => data_transfer_6_30_port, 
                           data_transfer(29) => data_transfer_6_29_port, 
                           data_transfer(28) => data_transfer_6_28_port, 
                           data_transfer(27) => data_transfer_6_27_port, 
                           data_transfer(26) => data_transfer_6_26_port, 
                           data_transfer(25) => data_transfer_6_25_port, 
                           data_transfer(24) => data_transfer_6_24_port, 
                           data_transfer(23) => data_transfer_6_23_port, 
                           data_transfer(22) => data_transfer_6_22_port, 
                           data_transfer(21) => data_transfer_6_21_port, 
                           data_transfer(20) => data_transfer_6_20_port, 
                           data_transfer(19) => data_transfer_6_19_port, 
                           data_transfer(18) => data_transfer_6_18_port, 
                           data_transfer(17) => data_transfer_6_17_port, 
                           data_transfer(16) => data_transfer_6_16_port, 
                           data_transfer(15) => data_transfer_6_15_port, 
                           data_transfer(14) => data_transfer_6_14_port, 
                           data_transfer(13) => data_transfer_6_13_port, 
                           data_transfer(12) => data_transfer_6_12_port, 
                           data_transfer(11) => data_transfer_6_11_port, 
                           data_transfer(10) => data_transfer_6_10_port, 
                           data_transfer(9) => data_transfer_6_9_port, 
                           data_transfer(8) => data_transfer_6_8_port, 
                           data_transfer(7) => data_transfer_6_7_port, 
                           data_transfer(6) => data_transfer_6_6_port, 
                           data_transfer(5) => data_transfer_6_5_port, 
                           data_transfer(4) => data_transfer_6_4_port, 
                           data_transfer(3) => data_transfer_6_3_port, 
                           data_transfer(2) => data_transfer_6_2_port, 
                           data_transfer(1) => data_transfer_6_1_port, 
                           data_transfer(0) => data_transfer_6_0_port, 
                           header(19) => header_12_PACKET_LENGTH_3_port, 
                           header(18) => header_12_PACKET_LENGTH_2_port, 
                           header(17) => header_12_PACKET_LENGTH_1_port, 
                           header(16) => header_12_PACKET_LENGTH_0_port, 
                           header(15) => header_12_X_DEST_1_port, header(14) =>
                           header_12_X_DEST_0_port, header(13) => 
                           header_12_Y_DEST_1_port, header(12) => 
                           header_12_Y_DEST_0_port, header(11) => 
                           header_12_Z_DEST_1_port, header(10) => 
                           header_12_Z_DEST_0_port, header(9) => 
                           header_11_PACKET_LENGTH_3_port, header(8) => 
                           header_11_PACKET_LENGTH_2_port, header(7) => 
                           header_11_PACKET_LENGTH_1_port, header(6) => 
                           header_11_PACKET_LENGTH_0_port, header(5) => 
                           header_11_X_DEST_1_port, header(4) => 
                           header_11_X_DEST_0_port, header(3) => 
                           header_11_Y_DEST_1_port, header(2) => 
                           header_11_Y_DEST_0_port, header(1) => 
                           header_11_Z_DEST_1_port, header(0) => 
                           header_11_Z_DEST_0_port);
   XBAR : crossbar_7_DXYU port map( crossbar_in(447) => data_transfer_6_63_port
                           , crossbar_in(446) => data_transfer_6_62_port, 
                           crossbar_in(445) => data_transfer_6_61_port, 
                           crossbar_in(444) => data_transfer_6_60_port, 
                           crossbar_in(443) => data_transfer_6_59_port, 
                           crossbar_in(442) => data_transfer_6_58_port, 
                           crossbar_in(441) => data_transfer_6_57_port, 
                           crossbar_in(440) => data_transfer_6_56_port, 
                           crossbar_in(439) => data_transfer_6_55_port, 
                           crossbar_in(438) => data_transfer_6_54_port, 
                           crossbar_in(437) => data_transfer_6_53_port, 
                           crossbar_in(436) => data_transfer_6_52_port, 
                           crossbar_in(435) => data_transfer_6_51_port, 
                           crossbar_in(434) => data_transfer_6_50_port, 
                           crossbar_in(433) => data_transfer_6_49_port, 
                           crossbar_in(432) => data_transfer_6_48_port, 
                           crossbar_in(431) => data_transfer_6_47_port, 
                           crossbar_in(430) => data_transfer_6_46_port, 
                           crossbar_in(429) => data_transfer_6_45_port, 
                           crossbar_in(428) => data_transfer_6_44_port, 
                           crossbar_in(427) => data_transfer_6_43_port, 
                           crossbar_in(426) => data_transfer_6_42_port, 
                           crossbar_in(425) => data_transfer_6_41_port, 
                           crossbar_in(424) => data_transfer_6_40_port, 
                           crossbar_in(423) => data_transfer_6_39_port, 
                           crossbar_in(422) => data_transfer_6_38_port, 
                           crossbar_in(421) => data_transfer_6_37_port, 
                           crossbar_in(420) => data_transfer_6_36_port, 
                           crossbar_in(419) => data_transfer_6_35_port, 
                           crossbar_in(418) => data_transfer_6_34_port, 
                           crossbar_in(417) => data_transfer_6_33_port, 
                           crossbar_in(416) => data_transfer_6_32_port, 
                           crossbar_in(415) => data_transfer_6_31_port, 
                           crossbar_in(414) => data_transfer_6_30_port, 
                           crossbar_in(413) => data_transfer_6_29_port, 
                           crossbar_in(412) => data_transfer_6_28_port, 
                           crossbar_in(411) => data_transfer_6_27_port, 
                           crossbar_in(410) => data_transfer_6_26_port, 
                           crossbar_in(409) => data_transfer_6_25_port, 
                           crossbar_in(408) => data_transfer_6_24_port, 
                           crossbar_in(407) => data_transfer_6_23_port, 
                           crossbar_in(406) => data_transfer_6_22_port, 
                           crossbar_in(405) => data_transfer_6_21_port, 
                           crossbar_in(404) => data_transfer_6_20_port, 
                           crossbar_in(403) => data_transfer_6_19_port, 
                           crossbar_in(402) => data_transfer_6_18_port, 
                           crossbar_in(401) => data_transfer_6_17_port, 
                           crossbar_in(400) => data_transfer_6_16_port, 
                           crossbar_in(399) => data_transfer_6_15_port, 
                           crossbar_in(398) => data_transfer_6_14_port, 
                           crossbar_in(397) => data_transfer_6_13_port, 
                           crossbar_in(396) => data_transfer_6_12_port, 
                           crossbar_in(395) => data_transfer_6_11_port, 
                           crossbar_in(394) => data_transfer_6_10_port, 
                           crossbar_in(393) => data_transfer_6_9_port, 
                           crossbar_in(392) => data_transfer_6_8_port, 
                           crossbar_in(391) => data_transfer_6_7_port, 
                           crossbar_in(390) => data_transfer_6_6_port, 
                           crossbar_in(389) => data_transfer_6_5_port, 
                           crossbar_in(388) => data_transfer_6_4_port, 
                           crossbar_in(387) => data_transfer_6_3_port, 
                           crossbar_in(386) => data_transfer_6_2_port, 
                           crossbar_in(385) => data_transfer_6_1_port, 
                           crossbar_in(384) => data_transfer_6_0_port, 
                           crossbar_in(383) => data_transfer_5_63_port, 
                           crossbar_in(382) => data_transfer_5_62_port, 
                           crossbar_in(381) => data_transfer_5_61_port, 
                           crossbar_in(380) => data_transfer_5_60_port, 
                           crossbar_in(379) => data_transfer_5_59_port, 
                           crossbar_in(378) => data_transfer_5_58_port, 
                           crossbar_in(377) => data_transfer_5_57_port, 
                           crossbar_in(376) => data_transfer_5_56_port, 
                           crossbar_in(375) => data_transfer_5_55_port, 
                           crossbar_in(374) => data_transfer_5_54_port, 
                           crossbar_in(373) => data_transfer_5_53_port, 
                           crossbar_in(372) => data_transfer_5_52_port, 
                           crossbar_in(371) => data_transfer_5_51_port, 
                           crossbar_in(370) => data_transfer_5_50_port, 
                           crossbar_in(369) => data_transfer_5_49_port, 
                           crossbar_in(368) => data_transfer_5_48_port, 
                           crossbar_in(367) => data_transfer_5_47_port, 
                           crossbar_in(366) => data_transfer_5_46_port, 
                           crossbar_in(365) => data_transfer_5_45_port, 
                           crossbar_in(364) => data_transfer_5_44_port, 
                           crossbar_in(363) => data_transfer_5_43_port, 
                           crossbar_in(362) => data_transfer_5_42_port, 
                           crossbar_in(361) => data_transfer_5_41_port, 
                           crossbar_in(360) => data_transfer_5_40_port, 
                           crossbar_in(359) => data_transfer_5_39_port, 
                           crossbar_in(358) => data_transfer_5_38_port, 
                           crossbar_in(357) => data_transfer_5_37_port, 
                           crossbar_in(356) => data_transfer_5_36_port, 
                           crossbar_in(355) => data_transfer_5_35_port, 
                           crossbar_in(354) => data_transfer_5_34_port, 
                           crossbar_in(353) => data_transfer_5_33_port, 
                           crossbar_in(352) => data_transfer_5_32_port, 
                           crossbar_in(351) => data_transfer_5_31_port, 
                           crossbar_in(350) => data_transfer_5_30_port, 
                           crossbar_in(349) => data_transfer_5_29_port, 
                           crossbar_in(348) => data_transfer_5_28_port, 
                           crossbar_in(347) => data_transfer_5_27_port, 
                           crossbar_in(346) => data_transfer_5_26_port, 
                           crossbar_in(345) => data_transfer_5_25_port, 
                           crossbar_in(344) => data_transfer_5_24_port, 
                           crossbar_in(343) => data_transfer_5_23_port, 
                           crossbar_in(342) => data_transfer_5_22_port, 
                           crossbar_in(341) => data_transfer_5_21_port, 
                           crossbar_in(340) => data_transfer_5_20_port, 
                           crossbar_in(339) => data_transfer_5_19_port, 
                           crossbar_in(338) => data_transfer_5_18_port, 
                           crossbar_in(337) => data_transfer_5_17_port, 
                           crossbar_in(336) => data_transfer_5_16_port, 
                           crossbar_in(335) => data_transfer_5_15_port, 
                           crossbar_in(334) => data_transfer_5_14_port, 
                           crossbar_in(333) => data_transfer_5_13_port, 
                           crossbar_in(332) => data_transfer_5_12_port, 
                           crossbar_in(331) => data_transfer_5_11_port, 
                           crossbar_in(330) => data_transfer_5_10_port, 
                           crossbar_in(329) => data_transfer_5_9_port, 
                           crossbar_in(328) => data_transfer_5_8_port, 
                           crossbar_in(327) => data_transfer_5_7_port, 
                           crossbar_in(326) => data_transfer_5_6_port, 
                           crossbar_in(325) => data_transfer_5_5_port, 
                           crossbar_in(324) => data_transfer_5_4_port, 
                           crossbar_in(323) => data_transfer_5_3_port, 
                           crossbar_in(322) => data_transfer_5_2_port, 
                           crossbar_in(321) => data_transfer_5_1_port, 
                           crossbar_in(320) => data_transfer_5_0_port, 
                           crossbar_in(319) => data_transfer_4_63_port, 
                           crossbar_in(318) => data_transfer_4_62_port, 
                           crossbar_in(317) => data_transfer_4_61_port, 
                           crossbar_in(316) => data_transfer_4_60_port, 
                           crossbar_in(315) => data_transfer_4_59_port, 
                           crossbar_in(314) => data_transfer_4_58_port, 
                           crossbar_in(313) => data_transfer_4_57_port, 
                           crossbar_in(312) => data_transfer_4_56_port, 
                           crossbar_in(311) => data_transfer_4_55_port, 
                           crossbar_in(310) => data_transfer_4_54_port, 
                           crossbar_in(309) => data_transfer_4_53_port, 
                           crossbar_in(308) => data_transfer_4_52_port, 
                           crossbar_in(307) => data_transfer_4_51_port, 
                           crossbar_in(306) => data_transfer_4_50_port, 
                           crossbar_in(305) => data_transfer_4_49_port, 
                           crossbar_in(304) => data_transfer_4_48_port, 
                           crossbar_in(303) => data_transfer_4_47_port, 
                           crossbar_in(302) => data_transfer_4_46_port, 
                           crossbar_in(301) => data_transfer_4_45_port, 
                           crossbar_in(300) => data_transfer_4_44_port, 
                           crossbar_in(299) => data_transfer_4_43_port, 
                           crossbar_in(298) => data_transfer_4_42_port, 
                           crossbar_in(297) => data_transfer_4_41_port, 
                           crossbar_in(296) => data_transfer_4_40_port, 
                           crossbar_in(295) => data_transfer_4_39_port, 
                           crossbar_in(294) => data_transfer_4_38_port, 
                           crossbar_in(293) => data_transfer_4_37_port, 
                           crossbar_in(292) => data_transfer_4_36_port, 
                           crossbar_in(291) => data_transfer_4_35_port, 
                           crossbar_in(290) => data_transfer_4_34_port, 
                           crossbar_in(289) => data_transfer_4_33_port, 
                           crossbar_in(288) => data_transfer_4_32_port, 
                           crossbar_in(287) => data_transfer_4_31_port, 
                           crossbar_in(286) => data_transfer_4_30_port, 
                           crossbar_in(285) => data_transfer_4_29_port, 
                           crossbar_in(284) => data_transfer_4_28_port, 
                           crossbar_in(283) => data_transfer_4_27_port, 
                           crossbar_in(282) => data_transfer_4_26_port, 
                           crossbar_in(281) => data_transfer_4_25_port, 
                           crossbar_in(280) => data_transfer_4_24_port, 
                           crossbar_in(279) => data_transfer_4_23_port, 
                           crossbar_in(278) => data_transfer_4_22_port, 
                           crossbar_in(277) => data_transfer_4_21_port, 
                           crossbar_in(276) => data_transfer_4_20_port, 
                           crossbar_in(275) => data_transfer_4_19_port, 
                           crossbar_in(274) => data_transfer_4_18_port, 
                           crossbar_in(273) => data_transfer_4_17_port, 
                           crossbar_in(272) => data_transfer_4_16_port, 
                           crossbar_in(271) => data_transfer_4_15_port, 
                           crossbar_in(270) => data_transfer_4_14_port, 
                           crossbar_in(269) => data_transfer_4_13_port, 
                           crossbar_in(268) => data_transfer_4_12_port, 
                           crossbar_in(267) => data_transfer_4_11_port, 
                           crossbar_in(266) => data_transfer_4_10_port, 
                           crossbar_in(265) => data_transfer_4_9_port, 
                           crossbar_in(264) => data_transfer_4_8_port, 
                           crossbar_in(263) => data_transfer_4_7_port, 
                           crossbar_in(262) => data_transfer_4_6_port, 
                           crossbar_in(261) => data_transfer_4_5_port, 
                           crossbar_in(260) => data_transfer_4_4_port, 
                           crossbar_in(259) => data_transfer_4_3_port, 
                           crossbar_in(258) => data_transfer_4_2_port, 
                           crossbar_in(257) => data_transfer_4_1_port, 
                           crossbar_in(256) => data_transfer_4_0_port, 
                           crossbar_in(255) => data_transfer_3_63_port, 
                           crossbar_in(254) => data_transfer_3_62_port, 
                           crossbar_in(253) => data_transfer_3_61_port, 
                           crossbar_in(252) => data_transfer_3_60_port, 
                           crossbar_in(251) => data_transfer_3_59_port, 
                           crossbar_in(250) => data_transfer_3_58_port, 
                           crossbar_in(249) => data_transfer_3_57_port, 
                           crossbar_in(248) => data_transfer_3_56_port, 
                           crossbar_in(247) => data_transfer_3_55_port, 
                           crossbar_in(246) => data_transfer_3_54_port, 
                           crossbar_in(245) => data_transfer_3_53_port, 
                           crossbar_in(244) => data_transfer_3_52_port, 
                           crossbar_in(243) => data_transfer_3_51_port, 
                           crossbar_in(242) => data_transfer_3_50_port, 
                           crossbar_in(241) => data_transfer_3_49_port, 
                           crossbar_in(240) => data_transfer_3_48_port, 
                           crossbar_in(239) => data_transfer_3_47_port, 
                           crossbar_in(238) => data_transfer_3_46_port, 
                           crossbar_in(237) => data_transfer_3_45_port, 
                           crossbar_in(236) => data_transfer_3_44_port, 
                           crossbar_in(235) => data_transfer_3_43_port, 
                           crossbar_in(234) => data_transfer_3_42_port, 
                           crossbar_in(233) => data_transfer_3_41_port, 
                           crossbar_in(232) => data_transfer_3_40_port, 
                           crossbar_in(231) => data_transfer_3_39_port, 
                           crossbar_in(230) => data_transfer_3_38_port, 
                           crossbar_in(229) => data_transfer_3_37_port, 
                           crossbar_in(228) => data_transfer_3_36_port, 
                           crossbar_in(227) => data_transfer_3_35_port, 
                           crossbar_in(226) => data_transfer_3_34_port, 
                           crossbar_in(225) => data_transfer_3_33_port, 
                           crossbar_in(224) => data_transfer_3_32_port, 
                           crossbar_in(223) => data_transfer_3_31_port, 
                           crossbar_in(222) => data_transfer_3_30_port, 
                           crossbar_in(221) => data_transfer_3_29_port, 
                           crossbar_in(220) => data_transfer_3_28_port, 
                           crossbar_in(219) => data_transfer_3_27_port, 
                           crossbar_in(218) => data_transfer_3_26_port, 
                           crossbar_in(217) => data_transfer_3_25_port, 
                           crossbar_in(216) => data_transfer_3_24_port, 
                           crossbar_in(215) => data_transfer_3_23_port, 
                           crossbar_in(214) => data_transfer_3_22_port, 
                           crossbar_in(213) => data_transfer_3_21_port, 
                           crossbar_in(212) => data_transfer_3_20_port, 
                           crossbar_in(211) => data_transfer_3_19_port, 
                           crossbar_in(210) => data_transfer_3_18_port, 
                           crossbar_in(209) => data_transfer_3_17_port, 
                           crossbar_in(208) => data_transfer_3_16_port, 
                           crossbar_in(207) => data_transfer_3_15_port, 
                           crossbar_in(206) => data_transfer_3_14_port, 
                           crossbar_in(205) => data_transfer_3_13_port, 
                           crossbar_in(204) => data_transfer_3_12_port, 
                           crossbar_in(203) => data_transfer_3_11_port, 
                           crossbar_in(202) => data_transfer_3_10_port, 
                           crossbar_in(201) => data_transfer_3_9_port, 
                           crossbar_in(200) => data_transfer_3_8_port, 
                           crossbar_in(199) => data_transfer_3_7_port, 
                           crossbar_in(198) => data_transfer_3_6_port, 
                           crossbar_in(197) => data_transfer_3_5_port, 
                           crossbar_in(196) => data_transfer_3_4_port, 
                           crossbar_in(195) => data_transfer_3_3_port, 
                           crossbar_in(194) => data_transfer_3_2_port, 
                           crossbar_in(193) => data_transfer_3_1_port, 
                           crossbar_in(192) => data_transfer_3_0_port, 
                           crossbar_in(191) => data_transfer_2_63_port, 
                           crossbar_in(190) => data_transfer_2_62_port, 
                           crossbar_in(189) => data_transfer_2_61_port, 
                           crossbar_in(188) => data_transfer_2_60_port, 
                           crossbar_in(187) => data_transfer_2_59_port, 
                           crossbar_in(186) => data_transfer_2_58_port, 
                           crossbar_in(185) => data_transfer_2_57_port, 
                           crossbar_in(184) => data_transfer_2_56_port, 
                           crossbar_in(183) => data_transfer_2_55_port, 
                           crossbar_in(182) => data_transfer_2_54_port, 
                           crossbar_in(181) => data_transfer_2_53_port, 
                           crossbar_in(180) => data_transfer_2_52_port, 
                           crossbar_in(179) => data_transfer_2_51_port, 
                           crossbar_in(178) => data_transfer_2_50_port, 
                           crossbar_in(177) => data_transfer_2_49_port, 
                           crossbar_in(176) => data_transfer_2_48_port, 
                           crossbar_in(175) => data_transfer_2_47_port, 
                           crossbar_in(174) => data_transfer_2_46_port, 
                           crossbar_in(173) => data_transfer_2_45_port, 
                           crossbar_in(172) => data_transfer_2_44_port, 
                           crossbar_in(171) => data_transfer_2_43_port, 
                           crossbar_in(170) => data_transfer_2_42_port, 
                           crossbar_in(169) => data_transfer_2_41_port, 
                           crossbar_in(168) => data_transfer_2_40_port, 
                           crossbar_in(167) => data_transfer_2_39_port, 
                           crossbar_in(166) => data_transfer_2_38_port, 
                           crossbar_in(165) => data_transfer_2_37_port, 
                           crossbar_in(164) => data_transfer_2_36_port, 
                           crossbar_in(163) => data_transfer_2_35_port, 
                           crossbar_in(162) => data_transfer_2_34_port, 
                           crossbar_in(161) => data_transfer_2_33_port, 
                           crossbar_in(160) => data_transfer_2_32_port, 
                           crossbar_in(159) => data_transfer_2_31_port, 
                           crossbar_in(158) => data_transfer_2_30_port, 
                           crossbar_in(157) => data_transfer_2_29_port, 
                           crossbar_in(156) => data_transfer_2_28_port, 
                           crossbar_in(155) => data_transfer_2_27_port, 
                           crossbar_in(154) => data_transfer_2_26_port, 
                           crossbar_in(153) => data_transfer_2_25_port, 
                           crossbar_in(152) => data_transfer_2_24_port, 
                           crossbar_in(151) => data_transfer_2_23_port, 
                           crossbar_in(150) => data_transfer_2_22_port, 
                           crossbar_in(149) => data_transfer_2_21_port, 
                           crossbar_in(148) => data_transfer_2_20_port, 
                           crossbar_in(147) => data_transfer_2_19_port, 
                           crossbar_in(146) => data_transfer_2_18_port, 
                           crossbar_in(145) => data_transfer_2_17_port, 
                           crossbar_in(144) => data_transfer_2_16_port, 
                           crossbar_in(143) => data_transfer_2_15_port, 
                           crossbar_in(142) => data_transfer_2_14_port, 
                           crossbar_in(141) => data_transfer_2_13_port, 
                           crossbar_in(140) => data_transfer_2_12_port, 
                           crossbar_in(139) => data_transfer_2_11_port, 
                           crossbar_in(138) => data_transfer_2_10_port, 
                           crossbar_in(137) => data_transfer_2_9_port, 
                           crossbar_in(136) => data_transfer_2_8_port, 
                           crossbar_in(135) => data_transfer_2_7_port, 
                           crossbar_in(134) => data_transfer_2_6_port, 
                           crossbar_in(133) => data_transfer_2_5_port, 
                           crossbar_in(132) => data_transfer_2_4_port, 
                           crossbar_in(131) => data_transfer_2_3_port, 
                           crossbar_in(130) => data_transfer_2_2_port, 
                           crossbar_in(129) => data_transfer_2_1_port, 
                           crossbar_in(128) => data_transfer_2_0_port, 
                           crossbar_in(127) => data_transfer_1_63_port, 
                           crossbar_in(126) => data_transfer_1_62_port, 
                           crossbar_in(125) => data_transfer_1_61_port, 
                           crossbar_in(124) => data_transfer_1_60_port, 
                           crossbar_in(123) => data_transfer_1_59_port, 
                           crossbar_in(122) => data_transfer_1_58_port, 
                           crossbar_in(121) => data_transfer_1_57_port, 
                           crossbar_in(120) => data_transfer_1_56_port, 
                           crossbar_in(119) => data_transfer_1_55_port, 
                           crossbar_in(118) => data_transfer_1_54_port, 
                           crossbar_in(117) => data_transfer_1_53_port, 
                           crossbar_in(116) => data_transfer_1_52_port, 
                           crossbar_in(115) => data_transfer_1_51_port, 
                           crossbar_in(114) => data_transfer_1_50_port, 
                           crossbar_in(113) => data_transfer_1_49_port, 
                           crossbar_in(112) => data_transfer_1_48_port, 
                           crossbar_in(111) => data_transfer_1_47_port, 
                           crossbar_in(110) => data_transfer_1_46_port, 
                           crossbar_in(109) => data_transfer_1_45_port, 
                           crossbar_in(108) => data_transfer_1_44_port, 
                           crossbar_in(107) => data_transfer_1_43_port, 
                           crossbar_in(106) => data_transfer_1_42_port, 
                           crossbar_in(105) => data_transfer_1_41_port, 
                           crossbar_in(104) => data_transfer_1_40_port, 
                           crossbar_in(103) => data_transfer_1_39_port, 
                           crossbar_in(102) => data_transfer_1_38_port, 
                           crossbar_in(101) => data_transfer_1_37_port, 
                           crossbar_in(100) => data_transfer_1_36_port, 
                           crossbar_in(99) => data_transfer_1_35_port, 
                           crossbar_in(98) => data_transfer_1_34_port, 
                           crossbar_in(97) => data_transfer_1_33_port, 
                           crossbar_in(96) => data_transfer_1_32_port, 
                           crossbar_in(95) => data_transfer_1_31_port, 
                           crossbar_in(94) => data_transfer_1_30_port, 
                           crossbar_in(93) => data_transfer_1_29_port, 
                           crossbar_in(92) => data_transfer_1_28_port, 
                           crossbar_in(91) => data_transfer_1_27_port, 
                           crossbar_in(90) => data_transfer_1_26_port, 
                           crossbar_in(89) => data_transfer_1_25_port, 
                           crossbar_in(88) => data_transfer_1_24_port, 
                           crossbar_in(87) => data_transfer_1_23_port, 
                           crossbar_in(86) => data_transfer_1_22_port, 
                           crossbar_in(85) => data_transfer_1_21_port, 
                           crossbar_in(84) => data_transfer_1_20_port, 
                           crossbar_in(83) => data_transfer_1_19_port, 
                           crossbar_in(82) => data_transfer_1_18_port, 
                           crossbar_in(81) => data_transfer_1_17_port, 
                           crossbar_in(80) => data_transfer_1_16_port, 
                           crossbar_in(79) => data_transfer_1_15_port, 
                           crossbar_in(78) => data_transfer_1_14_port, 
                           crossbar_in(77) => data_transfer_1_13_port, 
                           crossbar_in(76) => data_transfer_1_12_port, 
                           crossbar_in(75) => data_transfer_1_11_port, 
                           crossbar_in(74) => data_transfer_1_10_port, 
                           crossbar_in(73) => data_transfer_1_9_port, 
                           crossbar_in(72) => data_transfer_1_8_port, 
                           crossbar_in(71) => data_transfer_1_7_port, 
                           crossbar_in(70) => data_transfer_1_6_port, 
                           crossbar_in(69) => data_transfer_1_5_port, 
                           crossbar_in(68) => data_transfer_1_4_port, 
                           crossbar_in(67) => data_transfer_1_3_port, 
                           crossbar_in(66) => data_transfer_1_2_port, 
                           crossbar_in(65) => data_transfer_1_1_port, 
                           crossbar_in(64) => data_transfer_1_0_port, 
                           crossbar_in(63) => data_transfer_0_63_port, 
                           crossbar_in(62) => data_transfer_0_62_port, 
                           crossbar_in(61) => data_transfer_0_61_port, 
                           crossbar_in(60) => data_transfer_0_60_port, 
                           crossbar_in(59) => data_transfer_0_59_port, 
                           crossbar_in(58) => data_transfer_0_58_port, 
                           crossbar_in(57) => data_transfer_0_57_port, 
                           crossbar_in(56) => data_transfer_0_56_port, 
                           crossbar_in(55) => data_transfer_0_55_port, 
                           crossbar_in(54) => data_transfer_0_54_port, 
                           crossbar_in(53) => data_transfer_0_53_port, 
                           crossbar_in(52) => data_transfer_0_52_port, 
                           crossbar_in(51) => data_transfer_0_51_port, 
                           crossbar_in(50) => data_transfer_0_50_port, 
                           crossbar_in(49) => data_transfer_0_49_port, 
                           crossbar_in(48) => data_transfer_0_48_port, 
                           crossbar_in(47) => data_transfer_0_47_port, 
                           crossbar_in(46) => data_transfer_0_46_port, 
                           crossbar_in(45) => data_transfer_0_45_port, 
                           crossbar_in(44) => data_transfer_0_44_port, 
                           crossbar_in(43) => data_transfer_0_43_port, 
                           crossbar_in(42) => data_transfer_0_42_port, 
                           crossbar_in(41) => data_transfer_0_41_port, 
                           crossbar_in(40) => data_transfer_0_40_port, 
                           crossbar_in(39) => data_transfer_0_39_port, 
                           crossbar_in(38) => data_transfer_0_38_port, 
                           crossbar_in(37) => data_transfer_0_37_port, 
                           crossbar_in(36) => data_transfer_0_36_port, 
                           crossbar_in(35) => data_transfer_0_35_port, 
                           crossbar_in(34) => data_transfer_0_34_port, 
                           crossbar_in(33) => data_transfer_0_33_port, 
                           crossbar_in(32) => data_transfer_0_32_port, 
                           crossbar_in(31) => data_transfer_0_31_port, 
                           crossbar_in(30) => data_transfer_0_30_port, 
                           crossbar_in(29) => data_transfer_0_29_port, 
                           crossbar_in(28) => data_transfer_0_28_port, 
                           crossbar_in(27) => data_transfer_0_27_port, 
                           crossbar_in(26) => data_transfer_0_26_port, 
                           crossbar_in(25) => data_transfer_0_25_port, 
                           crossbar_in(24) => data_transfer_0_24_port, 
                           crossbar_in(23) => data_transfer_0_23_port, 
                           crossbar_in(22) => data_transfer_0_22_port, 
                           crossbar_in(21) => data_transfer_0_21_port, 
                           crossbar_in(20) => data_transfer_0_20_port, 
                           crossbar_in(19) => data_transfer_0_19_port, 
                           crossbar_in(18) => data_transfer_0_18_port, 
                           crossbar_in(17) => data_transfer_0_17_port, 
                           crossbar_in(16) => data_transfer_0_16_port, 
                           crossbar_in(15) => data_transfer_0_15_port, 
                           crossbar_in(14) => data_transfer_0_14_port, 
                           crossbar_in(13) => data_transfer_0_13_port, 
                           crossbar_in(12) => data_transfer_0_12_port, 
                           crossbar_in(11) => data_transfer_0_11_port, 
                           crossbar_in(10) => data_transfer_0_10_port, 
                           crossbar_in(9) => data_transfer_0_9_port, 
                           crossbar_in(8) => data_transfer_0_8_port, 
                           crossbar_in(7) => data_transfer_0_7_port, 
                           crossbar_in(6) => data_transfer_0_6_port, 
                           crossbar_in(5) => data_transfer_0_5_port, 
                           crossbar_in(4) => data_transfer_0_4_port, 
                           crossbar_in(3) => data_transfer_0_3_port, 
                           crossbar_in(2) => data_transfer_0_2_port, 
                           crossbar_in(1) => data_transfer_0_1_port, 
                           crossbar_in(0) => data_transfer_0_0_port, 
                           crossbar_ctrl(20) => crossbar_ctrl_20_port, 
                           crossbar_ctrl(19) => crossbar_ctrl_19_port, 
                           crossbar_ctrl(18) => crossbar_ctrl_18_port, 
                           crossbar_ctrl(17) => crossbar_ctrl_17_port, 
                           crossbar_ctrl(16) => crossbar_ctrl_16_port, 
                           crossbar_ctrl(15) => crossbar_ctrl_15_port, 
                           crossbar_ctrl(14) => crossbar_ctrl_14_port, 
                           crossbar_ctrl(13) => crossbar_ctrl_13_port, 
                           crossbar_ctrl(12) => crossbar_ctrl_12_port, 
                           crossbar_ctrl(11) => crossbar_ctrl_11_port, 
                           crossbar_ctrl(10) => crossbar_ctrl_10_port, 
                           crossbar_ctrl(9) => crossbar_ctrl_9_port, 
                           crossbar_ctrl(8) => crossbar_ctrl_8_port, 
                           crossbar_ctrl(7) => crossbar_ctrl_7_port, 
                           crossbar_ctrl(6) => crossbar_ctrl_6_port, 
                           crossbar_ctrl(5) => crossbar_ctrl_5_port, 
                           crossbar_ctrl(4) => crossbar_ctrl_4_port, 
                           crossbar_ctrl(3) => crossbar_ctrl_3_port, 
                           crossbar_ctrl(2) => crossbar_ctrl_2_port, 
                           crossbar_ctrl(1) => crossbar_ctrl_1_port, 
                           crossbar_ctrl(0) => crossbar_ctrl_0_port, 
                           crossbar_out(447) => data_tx_6_63_port, 
                           crossbar_out(446) => data_tx_6_62_port, 
                           crossbar_out(445) => data_tx_6_61_port, 
                           crossbar_out(444) => data_tx_6_60_port, 
                           crossbar_out(443) => data_tx_6_59_port, 
                           crossbar_out(442) => data_tx_6_58_port, 
                           crossbar_out(441) => data_tx_6_57_port, 
                           crossbar_out(440) => data_tx_6_56_port, 
                           crossbar_out(439) => data_tx_6_55_port, 
                           crossbar_out(438) => data_tx_6_54_port, 
                           crossbar_out(437) => data_tx_6_53_port, 
                           crossbar_out(436) => data_tx_6_52_port, 
                           crossbar_out(435) => data_tx_6_51_port, 
                           crossbar_out(434) => data_tx_6_50_port, 
                           crossbar_out(433) => data_tx_6_49_port, 
                           crossbar_out(432) => data_tx_6_48_port, 
                           crossbar_out(431) => data_tx_6_47_port, 
                           crossbar_out(430) => data_tx_6_46_port, 
                           crossbar_out(429) => data_tx_6_45_port, 
                           crossbar_out(428) => data_tx_6_44_port, 
                           crossbar_out(427) => data_tx_6_43_port, 
                           crossbar_out(426) => data_tx_6_42_port, 
                           crossbar_out(425) => data_tx_6_41_port, 
                           crossbar_out(424) => data_tx_6_40_port, 
                           crossbar_out(423) => data_tx_6_39_port, 
                           crossbar_out(422) => data_tx_6_38_port, 
                           crossbar_out(421) => data_tx_6_37_port, 
                           crossbar_out(420) => data_tx_6_36_port, 
                           crossbar_out(419) => data_tx_6_35_port, 
                           crossbar_out(418) => data_tx_6_34_port, 
                           crossbar_out(417) => data_tx_6_33_port, 
                           crossbar_out(416) => data_tx_6_32_port, 
                           crossbar_out(415) => data_tx_6_31_port, 
                           crossbar_out(414) => data_tx_6_30_port, 
                           crossbar_out(413) => data_tx_6_29_port, 
                           crossbar_out(412) => data_tx_6_28_port, 
                           crossbar_out(411) => data_tx_6_27_port, 
                           crossbar_out(410) => data_tx_6_26_port, 
                           crossbar_out(409) => data_tx_6_25_port, 
                           crossbar_out(408) => data_tx_6_24_port, 
                           crossbar_out(407) => data_tx_6_23_port, 
                           crossbar_out(406) => data_tx_6_22_port, 
                           crossbar_out(405) => data_tx_6_21_port, 
                           crossbar_out(404) => data_tx_6_20_port, 
                           crossbar_out(403) => data_tx_6_19_port, 
                           crossbar_out(402) => data_tx_6_18_port, 
                           crossbar_out(401) => data_tx_6_17_port, 
                           crossbar_out(400) => data_tx_6_16_port, 
                           crossbar_out(399) => data_tx_6_15_port, 
                           crossbar_out(398) => data_tx_6_14_port, 
                           crossbar_out(397) => data_tx_6_13_port, 
                           crossbar_out(396) => data_tx_6_12_port, 
                           crossbar_out(395) => data_tx_6_11_port, 
                           crossbar_out(394) => data_tx_6_10_port, 
                           crossbar_out(393) => data_tx_6_9_port, 
                           crossbar_out(392) => data_tx_6_8_port, 
                           crossbar_out(391) => data_tx_6_7_port, 
                           crossbar_out(390) => data_tx_6_6_port, 
                           crossbar_out(389) => data_tx_6_5_port, 
                           crossbar_out(388) => data_tx_6_4_port, 
                           crossbar_out(387) => data_tx_6_3_port, 
                           crossbar_out(386) => data_tx_6_2_port, 
                           crossbar_out(385) => data_tx_6_1_port, 
                           crossbar_out(384) => data_tx_6_0_port, 
                           crossbar_out(383) => data_tx_5_63_port, 
                           crossbar_out(382) => data_tx_5_62_port, 
                           crossbar_out(381) => data_tx_5_61_port, 
                           crossbar_out(380) => data_tx_5_60_port, 
                           crossbar_out(379) => data_tx_5_59_port, 
                           crossbar_out(378) => data_tx_5_58_port, 
                           crossbar_out(377) => data_tx_5_57_port, 
                           crossbar_out(376) => data_tx_5_56_port, 
                           crossbar_out(375) => data_tx_5_55_port, 
                           crossbar_out(374) => data_tx_5_54_port, 
                           crossbar_out(373) => data_tx_5_53_port, 
                           crossbar_out(372) => data_tx_5_52_port, 
                           crossbar_out(371) => data_tx_5_51_port, 
                           crossbar_out(370) => data_tx_5_50_port, 
                           crossbar_out(369) => data_tx_5_49_port, 
                           crossbar_out(368) => data_tx_5_48_port, 
                           crossbar_out(367) => data_tx_5_47_port, 
                           crossbar_out(366) => data_tx_5_46_port, 
                           crossbar_out(365) => data_tx_5_45_port, 
                           crossbar_out(364) => data_tx_5_44_port, 
                           crossbar_out(363) => data_tx_5_43_port, 
                           crossbar_out(362) => data_tx_5_42_port, 
                           crossbar_out(361) => data_tx_5_41_port, 
                           crossbar_out(360) => data_tx_5_40_port, 
                           crossbar_out(359) => data_tx_5_39_port, 
                           crossbar_out(358) => data_tx_5_38_port, 
                           crossbar_out(357) => data_tx_5_37_port, 
                           crossbar_out(356) => data_tx_5_36_port, 
                           crossbar_out(355) => data_tx_5_35_port, 
                           crossbar_out(354) => data_tx_5_34_port, 
                           crossbar_out(353) => data_tx_5_33_port, 
                           crossbar_out(352) => data_tx_5_32_port, 
                           crossbar_out(351) => data_tx_5_31_port, 
                           crossbar_out(350) => data_tx_5_30_port, 
                           crossbar_out(349) => data_tx_5_29_port, 
                           crossbar_out(348) => data_tx_5_28_port, 
                           crossbar_out(347) => data_tx_5_27_port, 
                           crossbar_out(346) => data_tx_5_26_port, 
                           crossbar_out(345) => data_tx_5_25_port, 
                           crossbar_out(344) => data_tx_5_24_port, 
                           crossbar_out(343) => data_tx_5_23_port, 
                           crossbar_out(342) => data_tx_5_22_port, 
                           crossbar_out(341) => data_tx_5_21_port, 
                           crossbar_out(340) => data_tx_5_20_port, 
                           crossbar_out(339) => data_tx_5_19_port, 
                           crossbar_out(338) => data_tx_5_18_port, 
                           crossbar_out(337) => data_tx_5_17_port, 
                           crossbar_out(336) => data_tx_5_16_port, 
                           crossbar_out(335) => data_tx_5_15_port, 
                           crossbar_out(334) => data_tx_5_14_port, 
                           crossbar_out(333) => data_tx_5_13_port, 
                           crossbar_out(332) => data_tx_5_12_port, 
                           crossbar_out(331) => data_tx_5_11_port, 
                           crossbar_out(330) => data_tx_5_10_port, 
                           crossbar_out(329) => data_tx_5_9_port, 
                           crossbar_out(328) => data_tx_5_8_port, 
                           crossbar_out(327) => data_tx_5_7_port, 
                           crossbar_out(326) => data_tx_5_6_port, 
                           crossbar_out(325) => data_tx_5_5_port, 
                           crossbar_out(324) => data_tx_5_4_port, 
                           crossbar_out(323) => data_tx_5_3_port, 
                           crossbar_out(322) => data_tx_5_2_port, 
                           crossbar_out(321) => data_tx_5_1_port, 
                           crossbar_out(320) => data_tx_5_0_port, 
                           crossbar_out(319) => data_tx_4_63_port, 
                           crossbar_out(318) => data_tx_4_62_port, 
                           crossbar_out(317) => data_tx_4_61_port, 
                           crossbar_out(316) => data_tx_4_60_port, 
                           crossbar_out(315) => data_tx_4_59_port, 
                           crossbar_out(314) => data_tx_4_58_port, 
                           crossbar_out(313) => data_tx_4_57_port, 
                           crossbar_out(312) => data_tx_4_56_port, 
                           crossbar_out(311) => data_tx_4_55_port, 
                           crossbar_out(310) => data_tx_4_54_port, 
                           crossbar_out(309) => data_tx_4_53_port, 
                           crossbar_out(308) => data_tx_4_52_port, 
                           crossbar_out(307) => data_tx_4_51_port, 
                           crossbar_out(306) => data_tx_4_50_port, 
                           crossbar_out(305) => data_tx_4_49_port, 
                           crossbar_out(304) => data_tx_4_48_port, 
                           crossbar_out(303) => data_tx_4_47_port, 
                           crossbar_out(302) => data_tx_4_46_port, 
                           crossbar_out(301) => data_tx_4_45_port, 
                           crossbar_out(300) => data_tx_4_44_port, 
                           crossbar_out(299) => data_tx_4_43_port, 
                           crossbar_out(298) => data_tx_4_42_port, 
                           crossbar_out(297) => data_tx_4_41_port, 
                           crossbar_out(296) => data_tx_4_40_port, 
                           crossbar_out(295) => data_tx_4_39_port, 
                           crossbar_out(294) => data_tx_4_38_port, 
                           crossbar_out(293) => data_tx_4_37_port, 
                           crossbar_out(292) => data_tx_4_36_port, 
                           crossbar_out(291) => data_tx_4_35_port, 
                           crossbar_out(290) => data_tx_4_34_port, 
                           crossbar_out(289) => data_tx_4_33_port, 
                           crossbar_out(288) => data_tx_4_32_port, 
                           crossbar_out(287) => data_tx_4_31_port, 
                           crossbar_out(286) => data_tx_4_30_port, 
                           crossbar_out(285) => data_tx_4_29_port, 
                           crossbar_out(284) => data_tx_4_28_port, 
                           crossbar_out(283) => data_tx_4_27_port, 
                           crossbar_out(282) => data_tx_4_26_port, 
                           crossbar_out(281) => data_tx_4_25_port, 
                           crossbar_out(280) => data_tx_4_24_port, 
                           crossbar_out(279) => data_tx_4_23_port, 
                           crossbar_out(278) => data_tx_4_22_port, 
                           crossbar_out(277) => data_tx_4_21_port, 
                           crossbar_out(276) => data_tx_4_20_port, 
                           crossbar_out(275) => data_tx_4_19_port, 
                           crossbar_out(274) => data_tx_4_18_port, 
                           crossbar_out(273) => data_tx_4_17_port, 
                           crossbar_out(272) => data_tx_4_16_port, 
                           crossbar_out(271) => data_tx_4_15_port, 
                           crossbar_out(270) => data_tx_4_14_port, 
                           crossbar_out(269) => data_tx_4_13_port, 
                           crossbar_out(268) => data_tx_4_12_port, 
                           crossbar_out(267) => data_tx_4_11_port, 
                           crossbar_out(266) => data_tx_4_10_port, 
                           crossbar_out(265) => data_tx_4_9_port, 
                           crossbar_out(264) => data_tx_4_8_port, 
                           crossbar_out(263) => data_tx_4_7_port, 
                           crossbar_out(262) => data_tx_4_6_port, 
                           crossbar_out(261) => data_tx_4_5_port, 
                           crossbar_out(260) => data_tx_4_4_port, 
                           crossbar_out(259) => data_tx_4_3_port, 
                           crossbar_out(258) => data_tx_4_2_port, 
                           crossbar_out(257) => data_tx_4_1_port, 
                           crossbar_out(256) => data_tx_4_0_port, 
                           crossbar_out(255) => data_tx_3_63_port, 
                           crossbar_out(254) => data_tx_3_62_port, 
                           crossbar_out(253) => data_tx_3_61_port, 
                           crossbar_out(252) => data_tx_3_60_port, 
                           crossbar_out(251) => data_tx_3_59_port, 
                           crossbar_out(250) => data_tx_3_58_port, 
                           crossbar_out(249) => data_tx_3_57_port, 
                           crossbar_out(248) => data_tx_3_56_port, 
                           crossbar_out(247) => data_tx_3_55_port, 
                           crossbar_out(246) => data_tx_3_54_port, 
                           crossbar_out(245) => data_tx_3_53_port, 
                           crossbar_out(244) => data_tx_3_52_port, 
                           crossbar_out(243) => data_tx_3_51_port, 
                           crossbar_out(242) => data_tx_3_50_port, 
                           crossbar_out(241) => data_tx_3_49_port, 
                           crossbar_out(240) => data_tx_3_48_port, 
                           crossbar_out(239) => data_tx_3_47_port, 
                           crossbar_out(238) => data_tx_3_46_port, 
                           crossbar_out(237) => data_tx_3_45_port, 
                           crossbar_out(236) => data_tx_3_44_port, 
                           crossbar_out(235) => data_tx_3_43_port, 
                           crossbar_out(234) => data_tx_3_42_port, 
                           crossbar_out(233) => data_tx_3_41_port, 
                           crossbar_out(232) => data_tx_3_40_port, 
                           crossbar_out(231) => data_tx_3_39_port, 
                           crossbar_out(230) => data_tx_3_38_port, 
                           crossbar_out(229) => data_tx_3_37_port, 
                           crossbar_out(228) => data_tx_3_36_port, 
                           crossbar_out(227) => data_tx_3_35_port, 
                           crossbar_out(226) => data_tx_3_34_port, 
                           crossbar_out(225) => data_tx_3_33_port, 
                           crossbar_out(224) => data_tx_3_32_port, 
                           crossbar_out(223) => data_tx_3_31_port, 
                           crossbar_out(222) => data_tx_3_30_port, 
                           crossbar_out(221) => data_tx_3_29_port, 
                           crossbar_out(220) => data_tx_3_28_port, 
                           crossbar_out(219) => data_tx_3_27_port, 
                           crossbar_out(218) => data_tx_3_26_port, 
                           crossbar_out(217) => data_tx_3_25_port, 
                           crossbar_out(216) => data_tx_3_24_port, 
                           crossbar_out(215) => data_tx_3_23_port, 
                           crossbar_out(214) => data_tx_3_22_port, 
                           crossbar_out(213) => data_tx_3_21_port, 
                           crossbar_out(212) => data_tx_3_20_port, 
                           crossbar_out(211) => data_tx_3_19_port, 
                           crossbar_out(210) => data_tx_3_18_port, 
                           crossbar_out(209) => data_tx_3_17_port, 
                           crossbar_out(208) => data_tx_3_16_port, 
                           crossbar_out(207) => data_tx_3_15_port, 
                           crossbar_out(206) => data_tx_3_14_port, 
                           crossbar_out(205) => data_tx_3_13_port, 
                           crossbar_out(204) => data_tx_3_12_port, 
                           crossbar_out(203) => data_tx_3_11_port, 
                           crossbar_out(202) => data_tx_3_10_port, 
                           crossbar_out(201) => data_tx_3_9_port, 
                           crossbar_out(200) => data_tx_3_8_port, 
                           crossbar_out(199) => data_tx_3_7_port, 
                           crossbar_out(198) => data_tx_3_6_port, 
                           crossbar_out(197) => data_tx_3_5_port, 
                           crossbar_out(196) => data_tx_3_4_port, 
                           crossbar_out(195) => data_tx_3_3_port, 
                           crossbar_out(194) => data_tx_3_2_port, 
                           crossbar_out(193) => data_tx_3_1_port, 
                           crossbar_out(192) => data_tx_3_0_port, 
                           crossbar_out(191) => data_tx_2_63_port, 
                           crossbar_out(190) => data_tx_2_62_port, 
                           crossbar_out(189) => data_tx_2_61_port, 
                           crossbar_out(188) => data_tx_2_60_port, 
                           crossbar_out(187) => data_tx_2_59_port, 
                           crossbar_out(186) => data_tx_2_58_port, 
                           crossbar_out(185) => data_tx_2_57_port, 
                           crossbar_out(184) => data_tx_2_56_port, 
                           crossbar_out(183) => data_tx_2_55_port, 
                           crossbar_out(182) => data_tx_2_54_port, 
                           crossbar_out(181) => data_tx_2_53_port, 
                           crossbar_out(180) => data_tx_2_52_port, 
                           crossbar_out(179) => data_tx_2_51_port, 
                           crossbar_out(178) => data_tx_2_50_port, 
                           crossbar_out(177) => data_tx_2_49_port, 
                           crossbar_out(176) => data_tx_2_48_port, 
                           crossbar_out(175) => data_tx_2_47_port, 
                           crossbar_out(174) => data_tx_2_46_port, 
                           crossbar_out(173) => data_tx_2_45_port, 
                           crossbar_out(172) => data_tx_2_44_port, 
                           crossbar_out(171) => data_tx_2_43_port, 
                           crossbar_out(170) => data_tx_2_42_port, 
                           crossbar_out(169) => data_tx_2_41_port, 
                           crossbar_out(168) => data_tx_2_40_port, 
                           crossbar_out(167) => data_tx_2_39_port, 
                           crossbar_out(166) => data_tx_2_38_port, 
                           crossbar_out(165) => data_tx_2_37_port, 
                           crossbar_out(164) => data_tx_2_36_port, 
                           crossbar_out(163) => data_tx_2_35_port, 
                           crossbar_out(162) => data_tx_2_34_port, 
                           crossbar_out(161) => data_tx_2_33_port, 
                           crossbar_out(160) => data_tx_2_32_port, 
                           crossbar_out(159) => data_tx_2_31_port, 
                           crossbar_out(158) => data_tx_2_30_port, 
                           crossbar_out(157) => data_tx_2_29_port, 
                           crossbar_out(156) => data_tx_2_28_port, 
                           crossbar_out(155) => data_tx_2_27_port, 
                           crossbar_out(154) => data_tx_2_26_port, 
                           crossbar_out(153) => data_tx_2_25_port, 
                           crossbar_out(152) => data_tx_2_24_port, 
                           crossbar_out(151) => data_tx_2_23_port, 
                           crossbar_out(150) => data_tx_2_22_port, 
                           crossbar_out(149) => data_tx_2_21_port, 
                           crossbar_out(148) => data_tx_2_20_port, 
                           crossbar_out(147) => data_tx_2_19_port, 
                           crossbar_out(146) => data_tx_2_18_port, 
                           crossbar_out(145) => data_tx_2_17_port, 
                           crossbar_out(144) => data_tx_2_16_port, 
                           crossbar_out(143) => data_tx_2_15_port, 
                           crossbar_out(142) => data_tx_2_14_port, 
                           crossbar_out(141) => data_tx_2_13_port, 
                           crossbar_out(140) => data_tx_2_12_port, 
                           crossbar_out(139) => data_tx_2_11_port, 
                           crossbar_out(138) => data_tx_2_10_port, 
                           crossbar_out(137) => data_tx_2_9_port, 
                           crossbar_out(136) => data_tx_2_8_port, 
                           crossbar_out(135) => data_tx_2_7_port, 
                           crossbar_out(134) => data_tx_2_6_port, 
                           crossbar_out(133) => data_tx_2_5_port, 
                           crossbar_out(132) => data_tx_2_4_port, 
                           crossbar_out(131) => data_tx_2_3_port, 
                           crossbar_out(130) => data_tx_2_2_port, 
                           crossbar_out(129) => data_tx_2_1_port, 
                           crossbar_out(128) => data_tx_2_0_port, 
                           crossbar_out(127) => data_tx_1_63_port, 
                           crossbar_out(126) => data_tx_1_62_port, 
                           crossbar_out(125) => data_tx_1_61_port, 
                           crossbar_out(124) => data_tx_1_60_port, 
                           crossbar_out(123) => data_tx_1_59_port, 
                           crossbar_out(122) => data_tx_1_58_port, 
                           crossbar_out(121) => data_tx_1_57_port, 
                           crossbar_out(120) => data_tx_1_56_port, 
                           crossbar_out(119) => data_tx_1_55_port, 
                           crossbar_out(118) => data_tx_1_54_port, 
                           crossbar_out(117) => data_tx_1_53_port, 
                           crossbar_out(116) => data_tx_1_52_port, 
                           crossbar_out(115) => data_tx_1_51_port, 
                           crossbar_out(114) => data_tx_1_50_port, 
                           crossbar_out(113) => data_tx_1_49_port, 
                           crossbar_out(112) => data_tx_1_48_port, 
                           crossbar_out(111) => data_tx_1_47_port, 
                           crossbar_out(110) => data_tx_1_46_port, 
                           crossbar_out(109) => data_tx_1_45_port, 
                           crossbar_out(108) => data_tx_1_44_port, 
                           crossbar_out(107) => data_tx_1_43_port, 
                           crossbar_out(106) => data_tx_1_42_port, 
                           crossbar_out(105) => data_tx_1_41_port, 
                           crossbar_out(104) => data_tx_1_40_port, 
                           crossbar_out(103) => data_tx_1_39_port, 
                           crossbar_out(102) => data_tx_1_38_port, 
                           crossbar_out(101) => data_tx_1_37_port, 
                           crossbar_out(100) => data_tx_1_36_port, 
                           crossbar_out(99) => data_tx_1_35_port, 
                           crossbar_out(98) => data_tx_1_34_port, 
                           crossbar_out(97) => data_tx_1_33_port, 
                           crossbar_out(96) => data_tx_1_32_port, 
                           crossbar_out(95) => data_tx_1_31_port, 
                           crossbar_out(94) => data_tx_1_30_port, 
                           crossbar_out(93) => data_tx_1_29_port, 
                           crossbar_out(92) => data_tx_1_28_port, 
                           crossbar_out(91) => data_tx_1_27_port, 
                           crossbar_out(90) => data_tx_1_26_port, 
                           crossbar_out(89) => data_tx_1_25_port, 
                           crossbar_out(88) => data_tx_1_24_port, 
                           crossbar_out(87) => data_tx_1_23_port, 
                           crossbar_out(86) => data_tx_1_22_port, 
                           crossbar_out(85) => data_tx_1_21_port, 
                           crossbar_out(84) => data_tx_1_20_port, 
                           crossbar_out(83) => data_tx_1_19_port, 
                           crossbar_out(82) => data_tx_1_18_port, 
                           crossbar_out(81) => data_tx_1_17_port, 
                           crossbar_out(80) => data_tx_1_16_port, 
                           crossbar_out(79) => data_tx_1_15_port, 
                           crossbar_out(78) => data_tx_1_14_port, 
                           crossbar_out(77) => data_tx_1_13_port, 
                           crossbar_out(76) => data_tx_1_12_port, 
                           crossbar_out(75) => data_tx_1_11_port, 
                           crossbar_out(74) => data_tx_1_10_port, 
                           crossbar_out(73) => data_tx_1_9_port, 
                           crossbar_out(72) => data_tx_1_8_port, 
                           crossbar_out(71) => data_tx_1_7_port, 
                           crossbar_out(70) => data_tx_1_6_port, 
                           crossbar_out(69) => data_tx_1_5_port, 
                           crossbar_out(68) => data_tx_1_4_port, 
                           crossbar_out(67) => data_tx_1_3_port, 
                           crossbar_out(66) => data_tx_1_2_port, 
                           crossbar_out(65) => data_tx_1_1_port, 
                           crossbar_out(64) => data_tx_1_0_port, 
                           crossbar_out(63) => data_tx_0_63_port, 
                           crossbar_out(62) => data_tx_0_62_port, 
                           crossbar_out(61) => data_tx_0_61_port, 
                           crossbar_out(60) => data_tx_0_60_port, 
                           crossbar_out(59) => data_tx_0_59_port, 
                           crossbar_out(58) => data_tx_0_58_port, 
                           crossbar_out(57) => data_tx_0_57_port, 
                           crossbar_out(56) => data_tx_0_56_port, 
                           crossbar_out(55) => data_tx_0_55_port, 
                           crossbar_out(54) => data_tx_0_54_port, 
                           crossbar_out(53) => data_tx_0_53_port, 
                           crossbar_out(52) => data_tx_0_52_port, 
                           crossbar_out(51) => data_tx_0_51_port, 
                           crossbar_out(50) => data_tx_0_50_port, 
                           crossbar_out(49) => data_tx_0_49_port, 
                           crossbar_out(48) => data_tx_0_48_port, 
                           crossbar_out(47) => data_tx_0_47_port, 
                           crossbar_out(46) => data_tx_0_46_port, 
                           crossbar_out(45) => data_tx_0_45_port, 
                           crossbar_out(44) => data_tx_0_44_port, 
                           crossbar_out(43) => data_tx_0_43_port, 
                           crossbar_out(42) => data_tx_0_42_port, 
                           crossbar_out(41) => data_tx_0_41_port, 
                           crossbar_out(40) => data_tx_0_40_port, 
                           crossbar_out(39) => data_tx_0_39_port, 
                           crossbar_out(38) => data_tx_0_38_port, 
                           crossbar_out(37) => data_tx_0_37_port, 
                           crossbar_out(36) => data_tx_0_36_port, 
                           crossbar_out(35) => data_tx_0_35_port, 
                           crossbar_out(34) => data_tx_0_34_port, 
                           crossbar_out(33) => data_tx_0_33_port, 
                           crossbar_out(32) => data_tx_0_32_port, 
                           crossbar_out(31) => data_tx_0_31_port, 
                           crossbar_out(30) => data_tx_0_30_port, 
                           crossbar_out(29) => data_tx_0_29_port, 
                           crossbar_out(28) => data_tx_0_28_port, 
                           crossbar_out(27) => data_tx_0_27_port, 
                           crossbar_out(26) => data_tx_0_26_port, 
                           crossbar_out(25) => data_tx_0_25_port, 
                           crossbar_out(24) => data_tx_0_24_port, 
                           crossbar_out(23) => data_tx_0_23_port, 
                           crossbar_out(22) => data_tx_0_22_port, 
                           crossbar_out(21) => data_tx_0_21_port, 
                           crossbar_out(20) => data_tx_0_20_port, 
                           crossbar_out(19) => data_tx_0_19_port, 
                           crossbar_out(18) => data_tx_0_18_port, 
                           crossbar_out(17) => data_tx_0_17_port, 
                           crossbar_out(16) => data_tx_0_16_port, 
                           crossbar_out(15) => data_tx_0_15_port, 
                           crossbar_out(14) => data_tx_0_14_port, 
                           crossbar_out(13) => data_tx_0_13_port, 
                           crossbar_out(12) => data_tx_0_12_port, 
                           crossbar_out(11) => data_tx_0_11_port, 
                           crossbar_out(10) => data_tx_0_10_port, 
                           crossbar_out(9) => data_tx_0_9_port, crossbar_out(8)
                           => data_tx_0_8_port, crossbar_out(7) => 
                           data_tx_0_7_port, crossbar_out(6) => 
                           data_tx_0_6_port, crossbar_out(5) => 
                           data_tx_0_5_port, crossbar_out(4) => 
                           data_tx_0_4_port, crossbar_out(3) => 
                           data_tx_0_3_port, crossbar_out(2) => 
                           data_tx_0_2_port, crossbar_out(1) => 
                           data_tx_0_1_port, crossbar_out(0) => 
                           data_tx_0_0_port);
   output_register_i_0 : output_register_vc_num1_vc_num_out1 port map( clk => 
                           clk, rst => rst, data_tx(63) => data_tx_0_63_port, 
                           data_tx(62) => data_tx_0_62_port, data_tx(61) => 
                           data_tx_0_61_port, data_tx(60) => data_tx_0_60_port,
                           data_tx(59) => data_tx_0_59_port, data_tx(58) => 
                           data_tx_0_58_port, data_tx(57) => data_tx_0_57_port,
                           data_tx(56) => data_tx_0_56_port, data_tx(55) => 
                           data_tx_0_55_port, data_tx(54) => data_tx_0_54_port,
                           data_tx(53) => data_tx_0_53_port, data_tx(52) => 
                           data_tx_0_52_port, data_tx(51) => data_tx_0_51_port,
                           data_tx(50) => data_tx_0_50_port, data_tx(49) => 
                           data_tx_0_49_port, data_tx(48) => data_tx_0_48_port,
                           data_tx(47) => data_tx_0_47_port, data_tx(46) => 
                           data_tx_0_46_port, data_tx(45) => data_tx_0_45_port,
                           data_tx(44) => data_tx_0_44_port, data_tx(43) => 
                           data_tx_0_43_port, data_tx(42) => data_tx_0_42_port,
                           data_tx(41) => data_tx_0_41_port, data_tx(40) => 
                           data_tx_0_40_port, data_tx(39) => data_tx_0_39_port,
                           data_tx(38) => data_tx_0_38_port, data_tx(37) => 
                           data_tx_0_37_port, data_tx(36) => data_tx_0_36_port,
                           data_tx(35) => data_tx_0_35_port, data_tx(34) => 
                           data_tx_0_34_port, data_tx(33) => data_tx_0_33_port,
                           data_tx(32) => data_tx_0_32_port, data_tx(31) => 
                           data_tx_0_31_port, data_tx(30) => data_tx_0_30_port,
                           data_tx(29) => data_tx_0_29_port, data_tx(28) => 
                           data_tx_0_28_port, data_tx(27) => data_tx_0_27_port,
                           data_tx(26) => data_tx_0_26_port, data_tx(25) => 
                           data_tx_0_25_port, data_tx(24) => data_tx_0_24_port,
                           data_tx(23) => data_tx_0_23_port, data_tx(22) => 
                           data_tx_0_22_port, data_tx(21) => data_tx_0_21_port,
                           data_tx(20) => data_tx_0_20_port, data_tx(19) => 
                           data_tx_0_19_port, data_tx(18) => data_tx_0_18_port,
                           data_tx(17) => data_tx_0_17_port, data_tx(16) => 
                           data_tx_0_16_port, data_tx(15) => data_tx_0_15_port,
                           data_tx(14) => data_tx_0_14_port, data_tx(13) => 
                           data_tx_0_13_port, data_tx(12) => data_tx_0_12_port,
                           data_tx(11) => data_tx_0_11_port, data_tx(10) => 
                           data_tx_0_10_port, data_tx(9) => data_tx_0_9_port, 
                           data_tx(8) => data_tx_0_8_port, data_tx(7) => 
                           data_tx_0_7_port, data_tx(6) => data_tx_0_6_port, 
                           data_tx(5) => data_tx_0_5_port, data_tx(4) => 
                           data_tx_0_4_port, data_tx(3) => data_tx_0_3_port, 
                           data_tx(2) => data_tx_0_2_port, data_tx(1) => 
                           data_tx_0_1_port, data_tx(0) => data_tx_0_0_port, 
                           vc_write_tx => vc_write_tx_vec_0_port, incr_tx => 
                           vc_transfer_vec_0_port, data_tx_pl(63) => 
                           data_tx_pl(0)(63), data_tx_pl(62) => 
                           data_tx_pl(0)(62), data_tx_pl(61) => 
                           data_tx_pl(0)(61), data_tx_pl(60) => 
                           data_tx_pl(0)(60), data_tx_pl(59) => 
                           data_tx_pl(0)(59), data_tx_pl(58) => 
                           data_tx_pl(0)(58), data_tx_pl(57) => 
                           data_tx_pl(0)(57), data_tx_pl(56) => 
                           data_tx_pl(0)(56), data_tx_pl(55) => 
                           data_tx_pl(0)(55), data_tx_pl(54) => 
                           data_tx_pl(0)(54), data_tx_pl(53) => 
                           data_tx_pl(0)(53), data_tx_pl(52) => 
                           data_tx_pl(0)(52), data_tx_pl(51) => 
                           data_tx_pl(0)(51), data_tx_pl(50) => 
                           data_tx_pl(0)(50), data_tx_pl(49) => 
                           data_tx_pl(0)(49), data_tx_pl(48) => 
                           data_tx_pl(0)(48), data_tx_pl(47) => 
                           data_tx_pl(0)(47), data_tx_pl(46) => 
                           data_tx_pl(0)(46), data_tx_pl(45) => 
                           data_tx_pl(0)(45), data_tx_pl(44) => 
                           data_tx_pl(0)(44), data_tx_pl(43) => 
                           data_tx_pl(0)(43), data_tx_pl(42) => 
                           data_tx_pl(0)(42), data_tx_pl(41) => 
                           data_tx_pl(0)(41), data_tx_pl(40) => 
                           data_tx_pl(0)(40), data_tx_pl(39) => 
                           data_tx_pl(0)(39), data_tx_pl(38) => 
                           data_tx_pl(0)(38), data_tx_pl(37) => 
                           data_tx_pl(0)(37), data_tx_pl(36) => 
                           data_tx_pl(0)(36), data_tx_pl(35) => 
                           data_tx_pl(0)(35), data_tx_pl(34) => 
                           data_tx_pl(0)(34), data_tx_pl(33) => 
                           data_tx_pl(0)(33), data_tx_pl(32) => 
                           data_tx_pl(0)(32), data_tx_pl(31) => 
                           data_tx_pl(0)(31), data_tx_pl(30) => 
                           data_tx_pl(0)(30), data_tx_pl(29) => 
                           data_tx_pl(0)(29), data_tx_pl(28) => 
                           data_tx_pl(0)(28), data_tx_pl(27) => 
                           data_tx_pl(0)(27), data_tx_pl(26) => 
                           data_tx_pl(0)(26), data_tx_pl(25) => 
                           data_tx_pl(0)(25), data_tx_pl(24) => 
                           data_tx_pl(0)(24), data_tx_pl(23) => 
                           data_tx_pl(0)(23), data_tx_pl(22) => 
                           data_tx_pl(0)(22), data_tx_pl(21) => 
                           data_tx_pl(0)(21), data_tx_pl(20) => 
                           data_tx_pl(0)(20), data_tx_pl(19) => 
                           data_tx_pl(0)(19), data_tx_pl(18) => 
                           data_tx_pl(0)(18), data_tx_pl(17) => 
                           data_tx_pl(0)(17), data_tx_pl(16) => 
                           data_tx_pl(0)(16), data_tx_pl(15) => 
                           data_tx_pl(0)(15), data_tx_pl(14) => 
                           data_tx_pl(0)(14), data_tx_pl(13) => 
                           data_tx_pl(0)(13), data_tx_pl(12) => 
                           data_tx_pl(0)(12), data_tx_pl(11) => 
                           data_tx_pl(0)(11), data_tx_pl(10) => 
                           data_tx_pl(0)(10), data_tx_pl(9) => data_tx_pl(0)(9)
                           , data_tx_pl(8) => data_tx_pl(0)(8), data_tx_pl(7) 
                           => data_tx_pl(0)(7), data_tx_pl(6) => 
                           data_tx_pl(0)(6), data_tx_pl(5) => data_tx_pl(0)(5),
                           data_tx_pl(4) => data_tx_pl(0)(4), data_tx_pl(3) => 
                           data_tx_pl(0)(3), data_tx_pl(2) => data_tx_pl(0)(2),
                           data_tx_pl(1) => data_tx_pl(0)(1), data_tx_pl(0) => 
                           data_tx_pl(0)(0), vc_write_tx_pl => 
                           vc_write_tx_pl_vec(0), incr_tx_pl => 
                           incr_tx_pl_vec(0));
   output_register_i_1 : output_register_vc_num2_vc_num_out2_0 port map( clk =>
                           clk, rst => rst, data_tx(63) => data_tx_1_63_port, 
                           data_tx(62) => data_tx_1_62_port, data_tx(61) => 
                           data_tx_1_61_port, data_tx(60) => data_tx_1_60_port,
                           data_tx(59) => data_tx_1_59_port, data_tx(58) => 
                           data_tx_1_58_port, data_tx(57) => data_tx_1_57_port,
                           data_tx(56) => data_tx_1_56_port, data_tx(55) => 
                           data_tx_1_55_port, data_tx(54) => data_tx_1_54_port,
                           data_tx(53) => data_tx_1_53_port, data_tx(52) => 
                           data_tx_1_52_port, data_tx(51) => data_tx_1_51_port,
                           data_tx(50) => data_tx_1_50_port, data_tx(49) => 
                           data_tx_1_49_port, data_tx(48) => data_tx_1_48_port,
                           data_tx(47) => data_tx_1_47_port, data_tx(46) => 
                           data_tx_1_46_port, data_tx(45) => data_tx_1_45_port,
                           data_tx(44) => data_tx_1_44_port, data_tx(43) => 
                           data_tx_1_43_port, data_tx(42) => data_tx_1_42_port,
                           data_tx(41) => data_tx_1_41_port, data_tx(40) => 
                           data_tx_1_40_port, data_tx(39) => data_tx_1_39_port,
                           data_tx(38) => data_tx_1_38_port, data_tx(37) => 
                           data_tx_1_37_port, data_tx(36) => data_tx_1_36_port,
                           data_tx(35) => data_tx_1_35_port, data_tx(34) => 
                           data_tx_1_34_port, data_tx(33) => data_tx_1_33_port,
                           data_tx(32) => data_tx_1_32_port, data_tx(31) => 
                           data_tx_1_31_port, data_tx(30) => data_tx_1_30_port,
                           data_tx(29) => data_tx_1_29_port, data_tx(28) => 
                           data_tx_1_28_port, data_tx(27) => data_tx_1_27_port,
                           data_tx(26) => data_tx_1_26_port, data_tx(25) => 
                           data_tx_1_25_port, data_tx(24) => data_tx_1_24_port,
                           data_tx(23) => data_tx_1_23_port, data_tx(22) => 
                           data_tx_1_22_port, data_tx(21) => data_tx_1_21_port,
                           data_tx(20) => data_tx_1_20_port, data_tx(19) => 
                           data_tx_1_19_port, data_tx(18) => data_tx_1_18_port,
                           data_tx(17) => data_tx_1_17_port, data_tx(16) => 
                           data_tx_1_16_port, data_tx(15) => data_tx_1_15_port,
                           data_tx(14) => data_tx_1_14_port, data_tx(13) => 
                           data_tx_1_13_port, data_tx(12) => data_tx_1_12_port,
                           data_tx(11) => data_tx_1_11_port, data_tx(10) => 
                           data_tx_1_10_port, data_tx(9) => data_tx_1_9_port, 
                           data_tx(8) => data_tx_1_8_port, data_tx(7) => 
                           data_tx_1_7_port, data_tx(6) => data_tx_1_6_port, 
                           data_tx(5) => data_tx_1_5_port, data_tx(4) => 
                           data_tx_1_4_port, data_tx(3) => data_tx_1_3_port, 
                           data_tx(2) => data_tx_1_2_port, data_tx(1) => 
                           data_tx_1_1_port, data_tx(0) => data_tx_1_0_port, 
                           vc_write_tx(1) => vc_write_tx_vec_2_port, 
                           vc_write_tx(0) => vc_write_tx_vec_1_port, incr_tx(1)
                           => vc_transfer_vec_2_port, incr_tx(0) => 
                           vc_transfer_vec_1_port, data_tx_pl(63) => 
                           data_tx_pl(1)(63), data_tx_pl(62) => 
                           data_tx_pl(1)(62), data_tx_pl(61) => 
                           data_tx_pl(1)(61), data_tx_pl(60) => 
                           data_tx_pl(1)(60), data_tx_pl(59) => 
                           data_tx_pl(1)(59), data_tx_pl(58) => 
                           data_tx_pl(1)(58), data_tx_pl(57) => 
                           data_tx_pl(1)(57), data_tx_pl(56) => 
                           data_tx_pl(1)(56), data_tx_pl(55) => 
                           data_tx_pl(1)(55), data_tx_pl(54) => 
                           data_tx_pl(1)(54), data_tx_pl(53) => 
                           data_tx_pl(1)(53), data_tx_pl(52) => 
                           data_tx_pl(1)(52), data_tx_pl(51) => 
                           data_tx_pl(1)(51), data_tx_pl(50) => 
                           data_tx_pl(1)(50), data_tx_pl(49) => 
                           data_tx_pl(1)(49), data_tx_pl(48) => 
                           data_tx_pl(1)(48), data_tx_pl(47) => 
                           data_tx_pl(1)(47), data_tx_pl(46) => 
                           data_tx_pl(1)(46), data_tx_pl(45) => 
                           data_tx_pl(1)(45), data_tx_pl(44) => 
                           data_tx_pl(1)(44), data_tx_pl(43) => 
                           data_tx_pl(1)(43), data_tx_pl(42) => 
                           data_tx_pl(1)(42), data_tx_pl(41) => 
                           data_tx_pl(1)(41), data_tx_pl(40) => 
                           data_tx_pl(1)(40), data_tx_pl(39) => 
                           data_tx_pl(1)(39), data_tx_pl(38) => 
                           data_tx_pl(1)(38), data_tx_pl(37) => 
                           data_tx_pl(1)(37), data_tx_pl(36) => 
                           data_tx_pl(1)(36), data_tx_pl(35) => 
                           data_tx_pl(1)(35), data_tx_pl(34) => 
                           data_tx_pl(1)(34), data_tx_pl(33) => 
                           data_tx_pl(1)(33), data_tx_pl(32) => 
                           data_tx_pl(1)(32), data_tx_pl(31) => 
                           data_tx_pl(1)(31), data_tx_pl(30) => 
                           data_tx_pl(1)(30), data_tx_pl(29) => 
                           data_tx_pl(1)(29), data_tx_pl(28) => 
                           data_tx_pl(1)(28), data_tx_pl(27) => 
                           data_tx_pl(1)(27), data_tx_pl(26) => 
                           data_tx_pl(1)(26), data_tx_pl(25) => 
                           data_tx_pl(1)(25), data_tx_pl(24) => 
                           data_tx_pl(1)(24), data_tx_pl(23) => 
                           data_tx_pl(1)(23), data_tx_pl(22) => 
                           data_tx_pl(1)(22), data_tx_pl(21) => 
                           data_tx_pl(1)(21), data_tx_pl(20) => 
                           data_tx_pl(1)(20), data_tx_pl(19) => 
                           data_tx_pl(1)(19), data_tx_pl(18) => 
                           data_tx_pl(1)(18), data_tx_pl(17) => 
                           data_tx_pl(1)(17), data_tx_pl(16) => 
                           data_tx_pl(1)(16), data_tx_pl(15) => 
                           data_tx_pl(1)(15), data_tx_pl(14) => 
                           data_tx_pl(1)(14), data_tx_pl(13) => 
                           data_tx_pl(1)(13), data_tx_pl(12) => 
                           data_tx_pl(1)(12), data_tx_pl(11) => 
                           data_tx_pl(1)(11), data_tx_pl(10) => 
                           data_tx_pl(1)(10), data_tx_pl(9) => data_tx_pl(1)(9)
                           , data_tx_pl(8) => data_tx_pl(1)(8), data_tx_pl(7) 
                           => data_tx_pl(1)(7), data_tx_pl(6) => 
                           data_tx_pl(1)(6), data_tx_pl(5) => data_tx_pl(1)(5),
                           data_tx_pl(4) => data_tx_pl(1)(4), data_tx_pl(3) => 
                           data_tx_pl(1)(3), data_tx_pl(2) => data_tx_pl(1)(2),
                           data_tx_pl(1) => data_tx_pl(1)(1), data_tx_pl(0) => 
                           data_tx_pl(1)(0), vc_write_tx_pl(1) => 
                           vc_write_tx_pl_vec(2), vc_write_tx_pl(0) => 
                           vc_write_tx_pl_vec(1), incr_tx_pl(1) => 
                           incr_tx_pl_vec(2), incr_tx_pl(0) => 
                           incr_tx_pl_vec(1));
   output_register_i_2 : output_register_vc_num2_vc_num_out2_5 port map( clk =>
                           clk, rst => rst, data_tx(63) => data_tx_2_63_port, 
                           data_tx(62) => data_tx_2_62_port, data_tx(61) => 
                           data_tx_2_61_port, data_tx(60) => data_tx_2_60_port,
                           data_tx(59) => data_tx_2_59_port, data_tx(58) => 
                           data_tx_2_58_port, data_tx(57) => data_tx_2_57_port,
                           data_tx(56) => data_tx_2_56_port, data_tx(55) => 
                           data_tx_2_55_port, data_tx(54) => data_tx_2_54_port,
                           data_tx(53) => data_tx_2_53_port, data_tx(52) => 
                           data_tx_2_52_port, data_tx(51) => data_tx_2_51_port,
                           data_tx(50) => data_tx_2_50_port, data_tx(49) => 
                           data_tx_2_49_port, data_tx(48) => data_tx_2_48_port,
                           data_tx(47) => data_tx_2_47_port, data_tx(46) => 
                           data_tx_2_46_port, data_tx(45) => data_tx_2_45_port,
                           data_tx(44) => data_tx_2_44_port, data_tx(43) => 
                           data_tx_2_43_port, data_tx(42) => data_tx_2_42_port,
                           data_tx(41) => data_tx_2_41_port, data_tx(40) => 
                           data_tx_2_40_port, data_tx(39) => data_tx_2_39_port,
                           data_tx(38) => data_tx_2_38_port, data_tx(37) => 
                           data_tx_2_37_port, data_tx(36) => data_tx_2_36_port,
                           data_tx(35) => data_tx_2_35_port, data_tx(34) => 
                           data_tx_2_34_port, data_tx(33) => data_tx_2_33_port,
                           data_tx(32) => data_tx_2_32_port, data_tx(31) => 
                           data_tx_2_31_port, data_tx(30) => data_tx_2_30_port,
                           data_tx(29) => data_tx_2_29_port, data_tx(28) => 
                           data_tx_2_28_port, data_tx(27) => data_tx_2_27_port,
                           data_tx(26) => data_tx_2_26_port, data_tx(25) => 
                           data_tx_2_25_port, data_tx(24) => data_tx_2_24_port,
                           data_tx(23) => data_tx_2_23_port, data_tx(22) => 
                           data_tx_2_22_port, data_tx(21) => data_tx_2_21_port,
                           data_tx(20) => data_tx_2_20_port, data_tx(19) => 
                           data_tx_2_19_port, data_tx(18) => data_tx_2_18_port,
                           data_tx(17) => data_tx_2_17_port, data_tx(16) => 
                           data_tx_2_16_port, data_tx(15) => data_tx_2_15_port,
                           data_tx(14) => data_tx_2_14_port, data_tx(13) => 
                           data_tx_2_13_port, data_tx(12) => data_tx_2_12_port,
                           data_tx(11) => data_tx_2_11_port, data_tx(10) => 
                           data_tx_2_10_port, data_tx(9) => data_tx_2_9_port, 
                           data_tx(8) => data_tx_2_8_port, data_tx(7) => 
                           data_tx_2_7_port, data_tx(6) => data_tx_2_6_port, 
                           data_tx(5) => data_tx_2_5_port, data_tx(4) => 
                           data_tx_2_4_port, data_tx(3) => data_tx_2_3_port, 
                           data_tx(2) => data_tx_2_2_port, data_tx(1) => 
                           data_tx_2_1_port, data_tx(0) => data_tx_2_0_port, 
                           vc_write_tx(1) => vc_write_tx_vec_4_port, 
                           vc_write_tx(0) => vc_write_tx_vec_3_port, incr_tx(1)
                           => vc_transfer_vec_4_port, incr_tx(0) => 
                           vc_transfer_vec_3_port, data_tx_pl(63) => 
                           data_tx_pl(2)(63), data_tx_pl(62) => 
                           data_tx_pl(2)(62), data_tx_pl(61) => 
                           data_tx_pl(2)(61), data_tx_pl(60) => 
                           data_tx_pl(2)(60), data_tx_pl(59) => 
                           data_tx_pl(2)(59), data_tx_pl(58) => 
                           data_tx_pl(2)(58), data_tx_pl(57) => 
                           data_tx_pl(2)(57), data_tx_pl(56) => 
                           data_tx_pl(2)(56), data_tx_pl(55) => 
                           data_tx_pl(2)(55), data_tx_pl(54) => 
                           data_tx_pl(2)(54), data_tx_pl(53) => 
                           data_tx_pl(2)(53), data_tx_pl(52) => 
                           data_tx_pl(2)(52), data_tx_pl(51) => 
                           data_tx_pl(2)(51), data_tx_pl(50) => 
                           data_tx_pl(2)(50), data_tx_pl(49) => 
                           data_tx_pl(2)(49), data_tx_pl(48) => 
                           data_tx_pl(2)(48), data_tx_pl(47) => 
                           data_tx_pl(2)(47), data_tx_pl(46) => 
                           data_tx_pl(2)(46), data_tx_pl(45) => 
                           data_tx_pl(2)(45), data_tx_pl(44) => 
                           data_tx_pl(2)(44), data_tx_pl(43) => 
                           data_tx_pl(2)(43), data_tx_pl(42) => 
                           data_tx_pl(2)(42), data_tx_pl(41) => 
                           data_tx_pl(2)(41), data_tx_pl(40) => 
                           data_tx_pl(2)(40), data_tx_pl(39) => 
                           data_tx_pl(2)(39), data_tx_pl(38) => 
                           data_tx_pl(2)(38), data_tx_pl(37) => 
                           data_tx_pl(2)(37), data_tx_pl(36) => 
                           data_tx_pl(2)(36), data_tx_pl(35) => 
                           data_tx_pl(2)(35), data_tx_pl(34) => 
                           data_tx_pl(2)(34), data_tx_pl(33) => 
                           data_tx_pl(2)(33), data_tx_pl(32) => 
                           data_tx_pl(2)(32), data_tx_pl(31) => 
                           data_tx_pl(2)(31), data_tx_pl(30) => 
                           data_tx_pl(2)(30), data_tx_pl(29) => 
                           data_tx_pl(2)(29), data_tx_pl(28) => 
                           data_tx_pl(2)(28), data_tx_pl(27) => 
                           data_tx_pl(2)(27), data_tx_pl(26) => 
                           data_tx_pl(2)(26), data_tx_pl(25) => 
                           data_tx_pl(2)(25), data_tx_pl(24) => 
                           data_tx_pl(2)(24), data_tx_pl(23) => 
                           data_tx_pl(2)(23), data_tx_pl(22) => 
                           data_tx_pl(2)(22), data_tx_pl(21) => 
                           data_tx_pl(2)(21), data_tx_pl(20) => 
                           data_tx_pl(2)(20), data_tx_pl(19) => 
                           data_tx_pl(2)(19), data_tx_pl(18) => 
                           data_tx_pl(2)(18), data_tx_pl(17) => 
                           data_tx_pl(2)(17), data_tx_pl(16) => 
                           data_tx_pl(2)(16), data_tx_pl(15) => 
                           data_tx_pl(2)(15), data_tx_pl(14) => 
                           data_tx_pl(2)(14), data_tx_pl(13) => 
                           data_tx_pl(2)(13), data_tx_pl(12) => 
                           data_tx_pl(2)(12), data_tx_pl(11) => 
                           data_tx_pl(2)(11), data_tx_pl(10) => 
                           data_tx_pl(2)(10), data_tx_pl(9) => data_tx_pl(2)(9)
                           , data_tx_pl(8) => data_tx_pl(2)(8), data_tx_pl(7) 
                           => data_tx_pl(2)(7), data_tx_pl(6) => 
                           data_tx_pl(2)(6), data_tx_pl(5) => data_tx_pl(2)(5),
                           data_tx_pl(4) => data_tx_pl(2)(4), data_tx_pl(3) => 
                           data_tx_pl(2)(3), data_tx_pl(2) => data_tx_pl(2)(2),
                           data_tx_pl(1) => data_tx_pl(2)(1), data_tx_pl(0) => 
                           data_tx_pl(2)(0), vc_write_tx_pl(1) => 
                           vc_write_tx_pl_vec(4), vc_write_tx_pl(0) => 
                           vc_write_tx_pl_vec(3), incr_tx_pl(1) => 
                           incr_tx_pl_vec(4), incr_tx_pl(0) => 
                           incr_tx_pl_vec(3));
   output_register_i_3 : output_register_vc_num2_vc_num_out2_4 port map( clk =>
                           clk, rst => rst, data_tx(63) => data_tx_3_63_port, 
                           data_tx(62) => data_tx_3_62_port, data_tx(61) => 
                           data_tx_3_61_port, data_tx(60) => data_tx_3_60_port,
                           data_tx(59) => data_tx_3_59_port, data_tx(58) => 
                           data_tx_3_58_port, data_tx(57) => data_tx_3_57_port,
                           data_tx(56) => data_tx_3_56_port, data_tx(55) => 
                           data_tx_3_55_port, data_tx(54) => data_tx_3_54_port,
                           data_tx(53) => data_tx_3_53_port, data_tx(52) => 
                           data_tx_3_52_port, data_tx(51) => data_tx_3_51_port,
                           data_tx(50) => data_tx_3_50_port, data_tx(49) => 
                           data_tx_3_49_port, data_tx(48) => data_tx_3_48_port,
                           data_tx(47) => data_tx_3_47_port, data_tx(46) => 
                           data_tx_3_46_port, data_tx(45) => data_tx_3_45_port,
                           data_tx(44) => data_tx_3_44_port, data_tx(43) => 
                           data_tx_3_43_port, data_tx(42) => data_tx_3_42_port,
                           data_tx(41) => data_tx_3_41_port, data_tx(40) => 
                           data_tx_3_40_port, data_tx(39) => data_tx_3_39_port,
                           data_tx(38) => data_tx_3_38_port, data_tx(37) => 
                           data_tx_3_37_port, data_tx(36) => data_tx_3_36_port,
                           data_tx(35) => data_tx_3_35_port, data_tx(34) => 
                           data_tx_3_34_port, data_tx(33) => data_tx_3_33_port,
                           data_tx(32) => data_tx_3_32_port, data_tx(31) => 
                           data_tx_3_31_port, data_tx(30) => data_tx_3_30_port,
                           data_tx(29) => data_tx_3_29_port, data_tx(28) => 
                           data_tx_3_28_port, data_tx(27) => data_tx_3_27_port,
                           data_tx(26) => data_tx_3_26_port, data_tx(25) => 
                           data_tx_3_25_port, data_tx(24) => data_tx_3_24_port,
                           data_tx(23) => data_tx_3_23_port, data_tx(22) => 
                           data_tx_3_22_port, data_tx(21) => data_tx_3_21_port,
                           data_tx(20) => data_tx_3_20_port, data_tx(19) => 
                           data_tx_3_19_port, data_tx(18) => data_tx_3_18_port,
                           data_tx(17) => data_tx_3_17_port, data_tx(16) => 
                           data_tx_3_16_port, data_tx(15) => data_tx_3_15_port,
                           data_tx(14) => data_tx_3_14_port, data_tx(13) => 
                           data_tx_3_13_port, data_tx(12) => data_tx_3_12_port,
                           data_tx(11) => data_tx_3_11_port, data_tx(10) => 
                           data_tx_3_10_port, data_tx(9) => data_tx_3_9_port, 
                           data_tx(8) => data_tx_3_8_port, data_tx(7) => 
                           data_tx_3_7_port, data_tx(6) => data_tx_3_6_port, 
                           data_tx(5) => data_tx_3_5_port, data_tx(4) => 
                           data_tx_3_4_port, data_tx(3) => data_tx_3_3_port, 
                           data_tx(2) => data_tx_3_2_port, data_tx(1) => 
                           data_tx_3_1_port, data_tx(0) => data_tx_3_0_port, 
                           vc_write_tx(1) => vc_write_tx_vec_6_port, 
                           vc_write_tx(0) => vc_write_tx_vec_5_port, incr_tx(1)
                           => vc_transfer_vec_6_port, incr_tx(0) => 
                           vc_transfer_vec_5_port, data_tx_pl(63) => 
                           data_tx_pl(3)(63), data_tx_pl(62) => 
                           data_tx_pl(3)(62), data_tx_pl(61) => 
                           data_tx_pl(3)(61), data_tx_pl(60) => 
                           data_tx_pl(3)(60), data_tx_pl(59) => 
                           data_tx_pl(3)(59), data_tx_pl(58) => 
                           data_tx_pl(3)(58), data_tx_pl(57) => 
                           data_tx_pl(3)(57), data_tx_pl(56) => 
                           data_tx_pl(3)(56), data_tx_pl(55) => 
                           data_tx_pl(3)(55), data_tx_pl(54) => 
                           data_tx_pl(3)(54), data_tx_pl(53) => 
                           data_tx_pl(3)(53), data_tx_pl(52) => 
                           data_tx_pl(3)(52), data_tx_pl(51) => 
                           data_tx_pl(3)(51), data_tx_pl(50) => 
                           data_tx_pl(3)(50), data_tx_pl(49) => 
                           data_tx_pl(3)(49), data_tx_pl(48) => 
                           data_tx_pl(3)(48), data_tx_pl(47) => 
                           data_tx_pl(3)(47), data_tx_pl(46) => 
                           data_tx_pl(3)(46), data_tx_pl(45) => 
                           data_tx_pl(3)(45), data_tx_pl(44) => 
                           data_tx_pl(3)(44), data_tx_pl(43) => 
                           data_tx_pl(3)(43), data_tx_pl(42) => 
                           data_tx_pl(3)(42), data_tx_pl(41) => 
                           data_tx_pl(3)(41), data_tx_pl(40) => 
                           data_tx_pl(3)(40), data_tx_pl(39) => 
                           data_tx_pl(3)(39), data_tx_pl(38) => 
                           data_tx_pl(3)(38), data_tx_pl(37) => 
                           data_tx_pl(3)(37), data_tx_pl(36) => 
                           data_tx_pl(3)(36), data_tx_pl(35) => 
                           data_tx_pl(3)(35), data_tx_pl(34) => 
                           data_tx_pl(3)(34), data_tx_pl(33) => 
                           data_tx_pl(3)(33), data_tx_pl(32) => 
                           data_tx_pl(3)(32), data_tx_pl(31) => 
                           data_tx_pl(3)(31), data_tx_pl(30) => 
                           data_tx_pl(3)(30), data_tx_pl(29) => 
                           data_tx_pl(3)(29), data_tx_pl(28) => 
                           data_tx_pl(3)(28), data_tx_pl(27) => 
                           data_tx_pl(3)(27), data_tx_pl(26) => 
                           data_tx_pl(3)(26), data_tx_pl(25) => 
                           data_tx_pl(3)(25), data_tx_pl(24) => 
                           data_tx_pl(3)(24), data_tx_pl(23) => 
                           data_tx_pl(3)(23), data_tx_pl(22) => 
                           data_tx_pl(3)(22), data_tx_pl(21) => 
                           data_tx_pl(3)(21), data_tx_pl(20) => 
                           data_tx_pl(3)(20), data_tx_pl(19) => 
                           data_tx_pl(3)(19), data_tx_pl(18) => 
                           data_tx_pl(3)(18), data_tx_pl(17) => 
                           data_tx_pl(3)(17), data_tx_pl(16) => 
                           data_tx_pl(3)(16), data_tx_pl(15) => 
                           data_tx_pl(3)(15), data_tx_pl(14) => 
                           data_tx_pl(3)(14), data_tx_pl(13) => 
                           data_tx_pl(3)(13), data_tx_pl(12) => 
                           data_tx_pl(3)(12), data_tx_pl(11) => 
                           data_tx_pl(3)(11), data_tx_pl(10) => 
                           data_tx_pl(3)(10), data_tx_pl(9) => data_tx_pl(3)(9)
                           , data_tx_pl(8) => data_tx_pl(3)(8), data_tx_pl(7) 
                           => data_tx_pl(3)(7), data_tx_pl(6) => 
                           data_tx_pl(3)(6), data_tx_pl(5) => data_tx_pl(3)(5),
                           data_tx_pl(4) => data_tx_pl(3)(4), data_tx_pl(3) => 
                           data_tx_pl(3)(3), data_tx_pl(2) => data_tx_pl(3)(2),
                           data_tx_pl(1) => data_tx_pl(3)(1), data_tx_pl(0) => 
                           data_tx_pl(3)(0), vc_write_tx_pl(1) => 
                           vc_write_tx_pl_vec(6), vc_write_tx_pl(0) => 
                           vc_write_tx_pl_vec(5), incr_tx_pl(1) => 
                           incr_tx_pl_vec(6), incr_tx_pl(0) => 
                           incr_tx_pl_vec(5));
   output_register_i_4 : output_register_vc_num2_vc_num_out2_3 port map( clk =>
                           clk, rst => rst, data_tx(63) => data_tx_4_63_port, 
                           data_tx(62) => data_tx_4_62_port, data_tx(61) => 
                           data_tx_4_61_port, data_tx(60) => data_tx_4_60_port,
                           data_tx(59) => data_tx_4_59_port, data_tx(58) => 
                           data_tx_4_58_port, data_tx(57) => data_tx_4_57_port,
                           data_tx(56) => data_tx_4_56_port, data_tx(55) => 
                           data_tx_4_55_port, data_tx(54) => data_tx_4_54_port,
                           data_tx(53) => data_tx_4_53_port, data_tx(52) => 
                           data_tx_4_52_port, data_tx(51) => data_tx_4_51_port,
                           data_tx(50) => data_tx_4_50_port, data_tx(49) => 
                           data_tx_4_49_port, data_tx(48) => data_tx_4_48_port,
                           data_tx(47) => data_tx_4_47_port, data_tx(46) => 
                           data_tx_4_46_port, data_tx(45) => data_tx_4_45_port,
                           data_tx(44) => data_tx_4_44_port, data_tx(43) => 
                           data_tx_4_43_port, data_tx(42) => data_tx_4_42_port,
                           data_tx(41) => data_tx_4_41_port, data_tx(40) => 
                           data_tx_4_40_port, data_tx(39) => data_tx_4_39_port,
                           data_tx(38) => data_tx_4_38_port, data_tx(37) => 
                           data_tx_4_37_port, data_tx(36) => data_tx_4_36_port,
                           data_tx(35) => data_tx_4_35_port, data_tx(34) => 
                           data_tx_4_34_port, data_tx(33) => data_tx_4_33_port,
                           data_tx(32) => data_tx_4_32_port, data_tx(31) => 
                           data_tx_4_31_port, data_tx(30) => data_tx_4_30_port,
                           data_tx(29) => data_tx_4_29_port, data_tx(28) => 
                           data_tx_4_28_port, data_tx(27) => data_tx_4_27_port,
                           data_tx(26) => data_tx_4_26_port, data_tx(25) => 
                           data_tx_4_25_port, data_tx(24) => data_tx_4_24_port,
                           data_tx(23) => data_tx_4_23_port, data_tx(22) => 
                           data_tx_4_22_port, data_tx(21) => data_tx_4_21_port,
                           data_tx(20) => data_tx_4_20_port, data_tx(19) => 
                           data_tx_4_19_port, data_tx(18) => data_tx_4_18_port,
                           data_tx(17) => data_tx_4_17_port, data_tx(16) => 
                           data_tx_4_16_port, data_tx(15) => data_tx_4_15_port,
                           data_tx(14) => data_tx_4_14_port, data_tx(13) => 
                           data_tx_4_13_port, data_tx(12) => data_tx_4_12_port,
                           data_tx(11) => data_tx_4_11_port, data_tx(10) => 
                           data_tx_4_10_port, data_tx(9) => data_tx_4_9_port, 
                           data_tx(8) => data_tx_4_8_port, data_tx(7) => 
                           data_tx_4_7_port, data_tx(6) => data_tx_4_6_port, 
                           data_tx(5) => data_tx_4_5_port, data_tx(4) => 
                           data_tx_4_4_port, data_tx(3) => data_tx_4_3_port, 
                           data_tx(2) => data_tx_4_2_port, data_tx(1) => 
                           data_tx_4_1_port, data_tx(0) => data_tx_4_0_port, 
                           vc_write_tx(1) => vc_write_tx_vec_8_port, 
                           vc_write_tx(0) => vc_write_tx_vec_7_port, incr_tx(1)
                           => vc_transfer_vec_8_port, incr_tx(0) => 
                           vc_transfer_vec_7_port, data_tx_pl(63) => 
                           data_tx_pl(4)(63), data_tx_pl(62) => 
                           data_tx_pl(4)(62), data_tx_pl(61) => 
                           data_tx_pl(4)(61), data_tx_pl(60) => 
                           data_tx_pl(4)(60), data_tx_pl(59) => 
                           data_tx_pl(4)(59), data_tx_pl(58) => 
                           data_tx_pl(4)(58), data_tx_pl(57) => 
                           data_tx_pl(4)(57), data_tx_pl(56) => 
                           data_tx_pl(4)(56), data_tx_pl(55) => 
                           data_tx_pl(4)(55), data_tx_pl(54) => 
                           data_tx_pl(4)(54), data_tx_pl(53) => 
                           data_tx_pl(4)(53), data_tx_pl(52) => 
                           data_tx_pl(4)(52), data_tx_pl(51) => 
                           data_tx_pl(4)(51), data_tx_pl(50) => 
                           data_tx_pl(4)(50), data_tx_pl(49) => 
                           data_tx_pl(4)(49), data_tx_pl(48) => 
                           data_tx_pl(4)(48), data_tx_pl(47) => 
                           data_tx_pl(4)(47), data_tx_pl(46) => 
                           data_tx_pl(4)(46), data_tx_pl(45) => 
                           data_tx_pl(4)(45), data_tx_pl(44) => 
                           data_tx_pl(4)(44), data_tx_pl(43) => 
                           data_tx_pl(4)(43), data_tx_pl(42) => 
                           data_tx_pl(4)(42), data_tx_pl(41) => 
                           data_tx_pl(4)(41), data_tx_pl(40) => 
                           data_tx_pl(4)(40), data_tx_pl(39) => 
                           data_tx_pl(4)(39), data_tx_pl(38) => 
                           data_tx_pl(4)(38), data_tx_pl(37) => 
                           data_tx_pl(4)(37), data_tx_pl(36) => 
                           data_tx_pl(4)(36), data_tx_pl(35) => 
                           data_tx_pl(4)(35), data_tx_pl(34) => 
                           data_tx_pl(4)(34), data_tx_pl(33) => 
                           data_tx_pl(4)(33), data_tx_pl(32) => 
                           data_tx_pl(4)(32), data_tx_pl(31) => 
                           data_tx_pl(4)(31), data_tx_pl(30) => 
                           data_tx_pl(4)(30), data_tx_pl(29) => 
                           data_tx_pl(4)(29), data_tx_pl(28) => 
                           data_tx_pl(4)(28), data_tx_pl(27) => 
                           data_tx_pl(4)(27), data_tx_pl(26) => 
                           data_tx_pl(4)(26), data_tx_pl(25) => 
                           data_tx_pl(4)(25), data_tx_pl(24) => 
                           data_tx_pl(4)(24), data_tx_pl(23) => 
                           data_tx_pl(4)(23), data_tx_pl(22) => 
                           data_tx_pl(4)(22), data_tx_pl(21) => 
                           data_tx_pl(4)(21), data_tx_pl(20) => 
                           data_tx_pl(4)(20), data_tx_pl(19) => 
                           data_tx_pl(4)(19), data_tx_pl(18) => 
                           data_tx_pl(4)(18), data_tx_pl(17) => 
                           data_tx_pl(4)(17), data_tx_pl(16) => 
                           data_tx_pl(4)(16), data_tx_pl(15) => 
                           data_tx_pl(4)(15), data_tx_pl(14) => 
                           data_tx_pl(4)(14), data_tx_pl(13) => 
                           data_tx_pl(4)(13), data_tx_pl(12) => 
                           data_tx_pl(4)(12), data_tx_pl(11) => 
                           data_tx_pl(4)(11), data_tx_pl(10) => 
                           data_tx_pl(4)(10), data_tx_pl(9) => data_tx_pl(4)(9)
                           , data_tx_pl(8) => data_tx_pl(4)(8), data_tx_pl(7) 
                           => data_tx_pl(4)(7), data_tx_pl(6) => 
                           data_tx_pl(4)(6), data_tx_pl(5) => data_tx_pl(4)(5),
                           data_tx_pl(4) => data_tx_pl(4)(4), data_tx_pl(3) => 
                           data_tx_pl(4)(3), data_tx_pl(2) => data_tx_pl(4)(2),
                           data_tx_pl(1) => data_tx_pl(4)(1), data_tx_pl(0) => 
                           data_tx_pl(4)(0), vc_write_tx_pl(1) => 
                           vc_write_tx_pl_vec(8), vc_write_tx_pl(0) => 
                           vc_write_tx_pl_vec(7), incr_tx_pl(1) => 
                           incr_tx_pl_vec(8), incr_tx_pl(0) => 
                           incr_tx_pl_vec(7));
   output_register_i_5 : output_register_vc_num2_vc_num_out2_2 port map( clk =>
                           clk, rst => rst, data_tx(63) => data_tx_5_63_port, 
                           data_tx(62) => data_tx_5_62_port, data_tx(61) => 
                           data_tx_5_61_port, data_tx(60) => data_tx_5_60_port,
                           data_tx(59) => data_tx_5_59_port, data_tx(58) => 
                           data_tx_5_58_port, data_tx(57) => data_tx_5_57_port,
                           data_tx(56) => data_tx_5_56_port, data_tx(55) => 
                           data_tx_5_55_port, data_tx(54) => data_tx_5_54_port,
                           data_tx(53) => data_tx_5_53_port, data_tx(52) => 
                           data_tx_5_52_port, data_tx(51) => data_tx_5_51_port,
                           data_tx(50) => data_tx_5_50_port, data_tx(49) => 
                           data_tx_5_49_port, data_tx(48) => data_tx_5_48_port,
                           data_tx(47) => data_tx_5_47_port, data_tx(46) => 
                           data_tx_5_46_port, data_tx(45) => data_tx_5_45_port,
                           data_tx(44) => data_tx_5_44_port, data_tx(43) => 
                           data_tx_5_43_port, data_tx(42) => data_tx_5_42_port,
                           data_tx(41) => data_tx_5_41_port, data_tx(40) => 
                           data_tx_5_40_port, data_tx(39) => data_tx_5_39_port,
                           data_tx(38) => data_tx_5_38_port, data_tx(37) => 
                           data_tx_5_37_port, data_tx(36) => data_tx_5_36_port,
                           data_tx(35) => data_tx_5_35_port, data_tx(34) => 
                           data_tx_5_34_port, data_tx(33) => data_tx_5_33_port,
                           data_tx(32) => data_tx_5_32_port, data_tx(31) => 
                           data_tx_5_31_port, data_tx(30) => data_tx_5_30_port,
                           data_tx(29) => data_tx_5_29_port, data_tx(28) => 
                           data_tx_5_28_port, data_tx(27) => data_tx_5_27_port,
                           data_tx(26) => data_tx_5_26_port, data_tx(25) => 
                           data_tx_5_25_port, data_tx(24) => data_tx_5_24_port,
                           data_tx(23) => data_tx_5_23_port, data_tx(22) => 
                           data_tx_5_22_port, data_tx(21) => data_tx_5_21_port,
                           data_tx(20) => data_tx_5_20_port, data_tx(19) => 
                           data_tx_5_19_port, data_tx(18) => data_tx_5_18_port,
                           data_tx(17) => data_tx_5_17_port, data_tx(16) => 
                           data_tx_5_16_port, data_tx(15) => data_tx_5_15_port,
                           data_tx(14) => data_tx_5_14_port, data_tx(13) => 
                           data_tx_5_13_port, data_tx(12) => data_tx_5_12_port,
                           data_tx(11) => data_tx_5_11_port, data_tx(10) => 
                           data_tx_5_10_port, data_tx(9) => data_tx_5_9_port, 
                           data_tx(8) => data_tx_5_8_port, data_tx(7) => 
                           data_tx_5_7_port, data_tx(6) => data_tx_5_6_port, 
                           data_tx(5) => data_tx_5_5_port, data_tx(4) => 
                           data_tx_5_4_port, data_tx(3) => data_tx_5_3_port, 
                           data_tx(2) => data_tx_5_2_port, data_tx(1) => 
                           data_tx_5_1_port, data_tx(0) => data_tx_5_0_port, 
                           vc_write_tx(1) => vc_write_tx_vec_10_port, 
                           vc_write_tx(0) => vc_write_tx_vec_9_port, incr_tx(1)
                           => vc_transfer_vec_10_port, incr_tx(0) => 
                           vc_transfer_vec_9_port, data_tx_pl(63) => 
                           data_tx_pl(5)(63), data_tx_pl(62) => 
                           data_tx_pl(5)(62), data_tx_pl(61) => 
                           data_tx_pl(5)(61), data_tx_pl(60) => 
                           data_tx_pl(5)(60), data_tx_pl(59) => 
                           data_tx_pl(5)(59), data_tx_pl(58) => 
                           data_tx_pl(5)(58), data_tx_pl(57) => 
                           data_tx_pl(5)(57), data_tx_pl(56) => 
                           data_tx_pl(5)(56), data_tx_pl(55) => 
                           data_tx_pl(5)(55), data_tx_pl(54) => 
                           data_tx_pl(5)(54), data_tx_pl(53) => 
                           data_tx_pl(5)(53), data_tx_pl(52) => 
                           data_tx_pl(5)(52), data_tx_pl(51) => 
                           data_tx_pl(5)(51), data_tx_pl(50) => 
                           data_tx_pl(5)(50), data_tx_pl(49) => 
                           data_tx_pl(5)(49), data_tx_pl(48) => 
                           data_tx_pl(5)(48), data_tx_pl(47) => 
                           data_tx_pl(5)(47), data_tx_pl(46) => 
                           data_tx_pl(5)(46), data_tx_pl(45) => 
                           data_tx_pl(5)(45), data_tx_pl(44) => 
                           data_tx_pl(5)(44), data_tx_pl(43) => 
                           data_tx_pl(5)(43), data_tx_pl(42) => 
                           data_tx_pl(5)(42), data_tx_pl(41) => 
                           data_tx_pl(5)(41), data_tx_pl(40) => 
                           data_tx_pl(5)(40), data_tx_pl(39) => 
                           data_tx_pl(5)(39), data_tx_pl(38) => 
                           data_tx_pl(5)(38), data_tx_pl(37) => 
                           data_tx_pl(5)(37), data_tx_pl(36) => 
                           data_tx_pl(5)(36), data_tx_pl(35) => 
                           data_tx_pl(5)(35), data_tx_pl(34) => 
                           data_tx_pl(5)(34), data_tx_pl(33) => 
                           data_tx_pl(5)(33), data_tx_pl(32) => 
                           data_tx_pl(5)(32), data_tx_pl(31) => 
                           data_tx_pl(5)(31), data_tx_pl(30) => 
                           data_tx_pl(5)(30), data_tx_pl(29) => 
                           data_tx_pl(5)(29), data_tx_pl(28) => 
                           data_tx_pl(5)(28), data_tx_pl(27) => 
                           data_tx_pl(5)(27), data_tx_pl(26) => 
                           data_tx_pl(5)(26), data_tx_pl(25) => 
                           data_tx_pl(5)(25), data_tx_pl(24) => 
                           data_tx_pl(5)(24), data_tx_pl(23) => 
                           data_tx_pl(5)(23), data_tx_pl(22) => 
                           data_tx_pl(5)(22), data_tx_pl(21) => 
                           data_tx_pl(5)(21), data_tx_pl(20) => 
                           data_tx_pl(5)(20), data_tx_pl(19) => 
                           data_tx_pl(5)(19), data_tx_pl(18) => 
                           data_tx_pl(5)(18), data_tx_pl(17) => 
                           data_tx_pl(5)(17), data_tx_pl(16) => 
                           data_tx_pl(5)(16), data_tx_pl(15) => 
                           data_tx_pl(5)(15), data_tx_pl(14) => 
                           data_tx_pl(5)(14), data_tx_pl(13) => 
                           data_tx_pl(5)(13), data_tx_pl(12) => 
                           data_tx_pl(5)(12), data_tx_pl(11) => 
                           data_tx_pl(5)(11), data_tx_pl(10) => 
                           data_tx_pl(5)(10), data_tx_pl(9) => data_tx_pl(5)(9)
                           , data_tx_pl(8) => data_tx_pl(5)(8), data_tx_pl(7) 
                           => data_tx_pl(5)(7), data_tx_pl(6) => 
                           data_tx_pl(5)(6), data_tx_pl(5) => data_tx_pl(5)(5),
                           data_tx_pl(4) => data_tx_pl(5)(4), data_tx_pl(3) => 
                           data_tx_pl(5)(3), data_tx_pl(2) => data_tx_pl(5)(2),
                           data_tx_pl(1) => data_tx_pl(5)(1), data_tx_pl(0) => 
                           data_tx_pl(5)(0), vc_write_tx_pl(1) => 
                           vc_write_tx_pl_vec(10), vc_write_tx_pl(0) => 
                           vc_write_tx_pl_vec(9), incr_tx_pl(1) => 
                           incr_tx_pl_vec(10), incr_tx_pl(0) => 
                           incr_tx_pl_vec(9));
   output_register_i_6 : output_register_vc_num2_vc_num_out2_1 port map( clk =>
                           clk, rst => rst, data_tx(63) => data_tx_6_63_port, 
                           data_tx(62) => data_tx_6_62_port, data_tx(61) => 
                           data_tx_6_61_port, data_tx(60) => data_tx_6_60_port,
                           data_tx(59) => data_tx_6_59_port, data_tx(58) => 
                           data_tx_6_58_port, data_tx(57) => data_tx_6_57_port,
                           data_tx(56) => data_tx_6_56_port, data_tx(55) => 
                           data_tx_6_55_port, data_tx(54) => data_tx_6_54_port,
                           data_tx(53) => data_tx_6_53_port, data_tx(52) => 
                           data_tx_6_52_port, data_tx(51) => data_tx_6_51_port,
                           data_tx(50) => data_tx_6_50_port, data_tx(49) => 
                           data_tx_6_49_port, data_tx(48) => data_tx_6_48_port,
                           data_tx(47) => data_tx_6_47_port, data_tx(46) => 
                           data_tx_6_46_port, data_tx(45) => data_tx_6_45_port,
                           data_tx(44) => data_tx_6_44_port, data_tx(43) => 
                           data_tx_6_43_port, data_tx(42) => data_tx_6_42_port,
                           data_tx(41) => data_tx_6_41_port, data_tx(40) => 
                           data_tx_6_40_port, data_tx(39) => data_tx_6_39_port,
                           data_tx(38) => data_tx_6_38_port, data_tx(37) => 
                           data_tx_6_37_port, data_tx(36) => data_tx_6_36_port,
                           data_tx(35) => data_tx_6_35_port, data_tx(34) => 
                           data_tx_6_34_port, data_tx(33) => data_tx_6_33_port,
                           data_tx(32) => data_tx_6_32_port, data_tx(31) => 
                           data_tx_6_31_port, data_tx(30) => data_tx_6_30_port,
                           data_tx(29) => data_tx_6_29_port, data_tx(28) => 
                           data_tx_6_28_port, data_tx(27) => data_tx_6_27_port,
                           data_tx(26) => data_tx_6_26_port, data_tx(25) => 
                           data_tx_6_25_port, data_tx(24) => data_tx_6_24_port,
                           data_tx(23) => data_tx_6_23_port, data_tx(22) => 
                           data_tx_6_22_port, data_tx(21) => data_tx_6_21_port,
                           data_tx(20) => data_tx_6_20_port, data_tx(19) => 
                           data_tx_6_19_port, data_tx(18) => data_tx_6_18_port,
                           data_tx(17) => data_tx_6_17_port, data_tx(16) => 
                           data_tx_6_16_port, data_tx(15) => data_tx_6_15_port,
                           data_tx(14) => data_tx_6_14_port, data_tx(13) => 
                           data_tx_6_13_port, data_tx(12) => data_tx_6_12_port,
                           data_tx(11) => data_tx_6_11_port, data_tx(10) => 
                           data_tx_6_10_port, data_tx(9) => data_tx_6_9_port, 
                           data_tx(8) => data_tx_6_8_port, data_tx(7) => 
                           data_tx_6_7_port, data_tx(6) => data_tx_6_6_port, 
                           data_tx(5) => data_tx_6_5_port, data_tx(4) => 
                           data_tx_6_4_port, data_tx(3) => data_tx_6_3_port, 
                           data_tx(2) => data_tx_6_2_port, data_tx(1) => 
                           data_tx_6_1_port, data_tx(0) => data_tx_6_0_port, 
                           vc_write_tx(1) => vc_write_tx_vec_12_port, 
                           vc_write_tx(0) => vc_write_tx_vec_11_port, 
                           incr_tx(1) => vc_transfer_vec_12_port, incr_tx(0) =>
                           vc_transfer_vec_11_port, data_tx_pl(63) => 
                           data_tx_pl(6)(63), data_tx_pl(62) => 
                           data_tx_pl(6)(62), data_tx_pl(61) => 
                           data_tx_pl(6)(61), data_tx_pl(60) => 
                           data_tx_pl(6)(60), data_tx_pl(59) => 
                           data_tx_pl(6)(59), data_tx_pl(58) => 
                           data_tx_pl(6)(58), data_tx_pl(57) => 
                           data_tx_pl(6)(57), data_tx_pl(56) => 
                           data_tx_pl(6)(56), data_tx_pl(55) => 
                           data_tx_pl(6)(55), data_tx_pl(54) => 
                           data_tx_pl(6)(54), data_tx_pl(53) => 
                           data_tx_pl(6)(53), data_tx_pl(52) => 
                           data_tx_pl(6)(52), data_tx_pl(51) => 
                           data_tx_pl(6)(51), data_tx_pl(50) => 
                           data_tx_pl(6)(50), data_tx_pl(49) => 
                           data_tx_pl(6)(49), data_tx_pl(48) => 
                           data_tx_pl(6)(48), data_tx_pl(47) => 
                           data_tx_pl(6)(47), data_tx_pl(46) => 
                           data_tx_pl(6)(46), data_tx_pl(45) => 
                           data_tx_pl(6)(45), data_tx_pl(44) => 
                           data_tx_pl(6)(44), data_tx_pl(43) => 
                           data_tx_pl(6)(43), data_tx_pl(42) => 
                           data_tx_pl(6)(42), data_tx_pl(41) => 
                           data_tx_pl(6)(41), data_tx_pl(40) => 
                           data_tx_pl(6)(40), data_tx_pl(39) => 
                           data_tx_pl(6)(39), data_tx_pl(38) => 
                           data_tx_pl(6)(38), data_tx_pl(37) => 
                           data_tx_pl(6)(37), data_tx_pl(36) => 
                           data_tx_pl(6)(36), data_tx_pl(35) => 
                           data_tx_pl(6)(35), data_tx_pl(34) => 
                           data_tx_pl(6)(34), data_tx_pl(33) => 
                           data_tx_pl(6)(33), data_tx_pl(32) => 
                           data_tx_pl(6)(32), data_tx_pl(31) => 
                           data_tx_pl(6)(31), data_tx_pl(30) => 
                           data_tx_pl(6)(30), data_tx_pl(29) => 
                           data_tx_pl(6)(29), data_tx_pl(28) => 
                           data_tx_pl(6)(28), data_tx_pl(27) => 
                           data_tx_pl(6)(27), data_tx_pl(26) => 
                           data_tx_pl(6)(26), data_tx_pl(25) => 
                           data_tx_pl(6)(25), data_tx_pl(24) => 
                           data_tx_pl(6)(24), data_tx_pl(23) => 
                           data_tx_pl(6)(23), data_tx_pl(22) => 
                           data_tx_pl(6)(22), data_tx_pl(21) => 
                           data_tx_pl(6)(21), data_tx_pl(20) => 
                           data_tx_pl(6)(20), data_tx_pl(19) => 
                           data_tx_pl(6)(19), data_tx_pl(18) => 
                           data_tx_pl(6)(18), data_tx_pl(17) => 
                           data_tx_pl(6)(17), data_tx_pl(16) => 
                           data_tx_pl(6)(16), data_tx_pl(15) => 
                           data_tx_pl(6)(15), data_tx_pl(14) => 
                           data_tx_pl(6)(14), data_tx_pl(13) => 
                           data_tx_pl(6)(13), data_tx_pl(12) => 
                           data_tx_pl(6)(12), data_tx_pl(11) => 
                           data_tx_pl(6)(11), data_tx_pl(10) => 
                           data_tx_pl(6)(10), data_tx_pl(9) => data_tx_pl(6)(9)
                           , data_tx_pl(8) => data_tx_pl(6)(8), data_tx_pl(7) 
                           => data_tx_pl(6)(7), data_tx_pl(6) => 
                           data_tx_pl(6)(6), data_tx_pl(5) => data_tx_pl(6)(5),
                           data_tx_pl(4) => data_tx_pl(6)(4), data_tx_pl(3) => 
                           data_tx_pl(6)(3), data_tx_pl(2) => data_tx_pl(6)(2),
                           data_tx_pl(1) => data_tx_pl(6)(1), data_tx_pl(0) => 
                           data_tx_pl(6)(0), vc_write_tx_pl(1) => 
                           vc_write_tx_pl_vec(12), vc_write_tx_pl(0) => 
                           vc_write_tx_pl_vec(11), incr_tx_pl(1) => 
                           incr_tx_pl_vec(12), incr_tx_pl(0) => 
                           incr_tx_pl_vec(11));
   CTRL_ARB : arbiter_7_1_1_1_1_DXYU port map( clk => clk, rst => rst, 
                           header(129) => header_12_PACKET_LENGTH_3_port, 
                           header(128) => header_12_PACKET_LENGTH_2_port, 
                           header(127) => header_12_PACKET_LENGTH_1_port, 
                           header(126) => header_12_PACKET_LENGTH_0_port, 
                           header(125) => header_12_X_DEST_1_port, header(124) 
                           => header_12_X_DEST_0_port, header(123) => 
                           header_12_Y_DEST_1_port, header(122) => 
                           header_12_Y_DEST_0_port, header(121) => 
                           header_12_Z_DEST_1_port, header(120) => 
                           header_12_Z_DEST_0_port, header(119) => 
                           header_11_PACKET_LENGTH_3_port, header(118) => 
                           header_11_PACKET_LENGTH_2_port, header(117) => 
                           header_11_PACKET_LENGTH_1_port, header(116) => 
                           header_11_PACKET_LENGTH_0_port, header(115) => 
                           header_11_X_DEST_1_port, header(114) => 
                           header_11_X_DEST_0_port, header(113) => 
                           header_11_Y_DEST_1_port, header(112) => 
                           header_11_Y_DEST_0_port, header(111) => 
                           header_11_Z_DEST_1_port, header(110) => 
                           header_11_Z_DEST_0_port, header(109) => 
                           header_10_PACKET_LENGTH_3_port, header(108) => 
                           header_10_PACKET_LENGTH_2_port, header(107) => 
                           header_10_PACKET_LENGTH_1_port, header(106) => 
                           header_10_PACKET_LENGTH_0_port, header(105) => 
                           header_10_X_DEST_1_port, header(104) => 
                           header_10_X_DEST_0_port, header(103) => 
                           header_10_Y_DEST_1_port, header(102) => 
                           header_10_Y_DEST_0_port, header(101) => 
                           header_10_Z_DEST_1_port, header(100) => 
                           header_10_Z_DEST_0_port, header(99) => 
                           header_9_PACKET_LENGTH_3_port, header(98) => 
                           header_9_PACKET_LENGTH_2_port, header(97) => 
                           header_9_PACKET_LENGTH_1_port, header(96) => 
                           header_9_PACKET_LENGTH_0_port, header(95) => 
                           header_9_X_DEST_1_port, header(94) => 
                           header_9_X_DEST_0_port, header(93) => 
                           header_9_Y_DEST_1_port, header(92) => 
                           header_9_Y_DEST_0_port, header(91) => 
                           header_9_Z_DEST_1_port, header(90) => 
                           header_9_Z_DEST_0_port, header(89) => 
                           header_8_PACKET_LENGTH_3_port, header(88) => 
                           header_8_PACKET_LENGTH_2_port, header(87) => 
                           header_8_PACKET_LENGTH_1_port, header(86) => 
                           header_8_PACKET_LENGTH_0_port, header(85) => 
                           header_8_X_DEST_1_port, header(84) => 
                           header_8_X_DEST_0_port, header(83) => 
                           header_8_Y_DEST_1_port, header(82) => 
                           header_8_Y_DEST_0_port, header(81) => 
                           header_8_Z_DEST_1_port, header(80) => 
                           header_8_Z_DEST_0_port, header(79) => 
                           header_7_PACKET_LENGTH_3_port, header(78) => 
                           header_7_PACKET_LENGTH_2_port, header(77) => 
                           header_7_PACKET_LENGTH_1_port, header(76) => 
                           header_7_PACKET_LENGTH_0_port, header(75) => 
                           header_7_X_DEST_1_port, header(74) => 
                           header_7_X_DEST_0_port, header(73) => 
                           header_7_Y_DEST_1_port, header(72) => 
                           header_7_Y_DEST_0_port, header(71) => 
                           header_7_Z_DEST_1_port, header(70) => 
                           header_7_Z_DEST_0_port, header(69) => 
                           header_6_PACKET_LENGTH_3_port, header(68) => 
                           header_6_PACKET_LENGTH_2_port, header(67) => 
                           header_6_PACKET_LENGTH_1_port, header(66) => 
                           header_6_PACKET_LENGTH_0_port, header(65) => 
                           header_6_X_DEST_1_port, header(64) => 
                           header_6_X_DEST_0_port, header(63) => 
                           header_6_Y_DEST_1_port, header(62) => 
                           header_6_Y_DEST_0_port, header(61) => 
                           header_6_Z_DEST_1_port, header(60) => 
                           header_6_Z_DEST_0_port, header(59) => 
                           header_5_PACKET_LENGTH_3_port, header(58) => 
                           header_5_PACKET_LENGTH_2_port, header(57) => 
                           header_5_PACKET_LENGTH_1_port, header(56) => 
                           header_5_PACKET_LENGTH_0_port, header(55) => 
                           header_5_X_DEST_1_port, header(54) => 
                           header_5_X_DEST_0_port, header(53) => 
                           header_5_Y_DEST_1_port, header(52) => 
                           header_5_Y_DEST_0_port, header(51) => 
                           header_5_Z_DEST_1_port, header(50) => 
                           header_5_Z_DEST_0_port, header(49) => 
                           header_4_PACKET_LENGTH_3_port, header(48) => 
                           header_4_PACKET_LENGTH_2_port, header(47) => 
                           header_4_PACKET_LENGTH_1_port, header(46) => 
                           header_4_PACKET_LENGTH_0_port, header(45) => 
                           header_4_X_DEST_1_port, header(44) => 
                           header_4_X_DEST_0_port, header(43) => 
                           header_4_Y_DEST_1_port, header(42) => 
                           header_4_Y_DEST_0_port, header(41) => 
                           header_4_Z_DEST_1_port, header(40) => 
                           header_4_Z_DEST_0_port, header(39) => 
                           header_3_PACKET_LENGTH_3_port, header(38) => 
                           header_3_PACKET_LENGTH_2_port, header(37) => 
                           header_3_PACKET_LENGTH_1_port, header(36) => 
                           header_3_PACKET_LENGTH_0_port, header(35) => 
                           header_3_X_DEST_1_port, header(34) => 
                           header_3_X_DEST_0_port, header(33) => 
                           header_3_Y_DEST_1_port, header(32) => 
                           header_3_Y_DEST_0_port, header(31) => 
                           header_3_Z_DEST_1_port, header(30) => 
                           header_3_Z_DEST_0_port, header(29) => 
                           header_2_PACKET_LENGTH_3_port, header(28) => 
                           header_2_PACKET_LENGTH_2_port, header(27) => 
                           header_2_PACKET_LENGTH_1_port, header(26) => 
                           header_2_PACKET_LENGTH_0_port, header(25) => 
                           header_2_X_DEST_1_port, header(24) => 
                           header_2_X_DEST_0_port, header(23) => 
                           header_2_Y_DEST_1_port, header(22) => 
                           header_2_Y_DEST_0_port, header(21) => 
                           header_2_Z_DEST_1_port, header(20) => 
                           header_2_Z_DEST_0_port, header(19) => 
                           header_1_PACKET_LENGTH_3_port, header(18) => 
                           header_1_PACKET_LENGTH_2_port, header(17) => 
                           header_1_PACKET_LENGTH_1_port, header(16) => 
                           header_1_PACKET_LENGTH_0_port, header(15) => 
                           header_1_X_DEST_1_port, header(14) => 
                           header_1_X_DEST_0_port, header(13) => 
                           header_1_Y_DEST_1_port, header(12) => 
                           header_1_Y_DEST_0_port, header(11) => 
                           header_1_Z_DEST_1_port, header(10) => 
                           header_1_Z_DEST_0_port, header(9) => 
                           header_0_PACKET_LENGTH_3_port, header(8) => 
                           header_0_PACKET_LENGTH_2_port, header(7) => 
                           header_0_PACKET_LENGTH_1_port, header(6) => 
                           header_0_PACKET_LENGTH_0_port, header(5) => 
                           header_0_X_DEST_1_port, header(4) => 
                           header_0_X_DEST_0_port, header(3) => 
                           header_0_Y_DEST_1_port, header(2) => 
                           header_0_Y_DEST_0_port, header(1) => 
                           header_0_Z_DEST_1_port, header(0) => 
                           header_0_Z_DEST_0_port, valid_data_vc_vec(12) => 
                           valid_data_vc_vec_12_port, valid_data_vc_vec(11) => 
                           valid_data_vc_vec_11_port, valid_data_vc_vec(10) => 
                           valid_data_vc_vec_10_port, valid_data_vc_vec(9) => 
                           valid_data_vc_vec_9_port, valid_data_vc_vec(8) => 
                           valid_data_vc_vec_8_port, valid_data_vc_vec(7) => 
                           valid_data_vc_vec_7_port, valid_data_vc_vec(6) => 
                           valid_data_vc_vec_6_port, valid_data_vc_vec(5) => 
                           valid_data_vc_vec_5_port, valid_data_vc_vec(4) => 
                           valid_data_vc_vec_4_port, valid_data_vc_vec(3) => 
                           valid_data_vc_vec_3_port, valid_data_vc_vec(2) => 
                           valid_data_vc_vec_2_port, valid_data_vc_vec(1) => 
                           valid_data_vc_vec_1_port, valid_data_vc_vec(0) => 
                           valid_data_vc_vec_0_port, incr_rx_vec(12) => 
                           incr_rx_vec(12), incr_rx_vec(11) => incr_rx_vec(11),
                           incr_rx_vec(10) => incr_rx_vec(10), incr_rx_vec(9) 
                           => incr_rx_vec(9), incr_rx_vec(8) => incr_rx_vec(8),
                           incr_rx_vec(7) => incr_rx_vec(7), incr_rx_vec(6) => 
                           incr_rx_vec(6), incr_rx_vec(5) => incr_rx_vec(5), 
                           incr_rx_vec(4) => incr_rx_vec(4), incr_rx_vec(3) => 
                           incr_rx_vec(3), incr_rx_vec(2) => incr_rx_vec(2), 
                           incr_rx_vec(1) => incr_rx_vec(1), incr_rx_vec(0) => 
                           incr_rx_vec(0), crossbar_ctrl(20) => 
                           crossbar_ctrl_20_port, crossbar_ctrl(19) => 
                           crossbar_ctrl_19_port, crossbar_ctrl(18) => 
                           crossbar_ctrl_18_port, crossbar_ctrl(17) => 
                           crossbar_ctrl_17_port, crossbar_ctrl(16) => 
                           crossbar_ctrl_16_port, crossbar_ctrl(15) => 
                           crossbar_ctrl_15_port, crossbar_ctrl(14) => 
                           crossbar_ctrl_14_port, crossbar_ctrl(13) => 
                           crossbar_ctrl_13_port, crossbar_ctrl(12) => 
                           crossbar_ctrl_12_port, crossbar_ctrl(11) => 
                           crossbar_ctrl_11_port, crossbar_ctrl(10) => 
                           crossbar_ctrl_10_port, crossbar_ctrl(9) => 
                           crossbar_ctrl_9_port, crossbar_ctrl(8) => 
                           crossbar_ctrl_8_port, crossbar_ctrl(7) => 
                           crossbar_ctrl_7_port, crossbar_ctrl(6) => 
                           crossbar_ctrl_6_port, crossbar_ctrl(5) => 
                           crossbar_ctrl_5_port, crossbar_ctrl(4) => 
                           crossbar_ctrl_4_port, crossbar_ctrl(3) => 
                           crossbar_ctrl_3_port, crossbar_ctrl(2) => 
                           crossbar_ctrl_2_port, crossbar_ctrl(1) => 
                           crossbar_ctrl_1_port, crossbar_ctrl(0) => 
                           crossbar_ctrl_0_port, vc_transfer_vec(12) => 
                           vc_transfer_vec_12_port, vc_transfer_vec(11) => 
                           vc_transfer_vec_11_port, vc_transfer_vec(10) => 
                           vc_transfer_vec_10_port, vc_transfer_vec(9) => 
                           vc_transfer_vec_9_port, vc_transfer_vec(8) => 
                           vc_transfer_vec_8_port, vc_transfer_vec(7) => 
                           vc_transfer_vec_7_port, vc_transfer_vec(6) => 
                           vc_transfer_vec_6_port, vc_transfer_vec(5) => 
                           vc_transfer_vec_5_port, vc_transfer_vec(4) => 
                           vc_transfer_vec_4_port, vc_transfer_vec(3) => 
                           vc_transfer_vec_3_port, vc_transfer_vec(2) => 
                           vc_transfer_vec_2_port, vc_transfer_vec(1) => 
                           vc_transfer_vec_1_port, vc_transfer_vec(0) => 
                           vc_transfer_vec_0_port, vc_write_tx_vec(12) => 
                           vc_write_tx_vec_12_port, vc_write_tx_vec(11) => 
                           vc_write_tx_vec_11_port, vc_write_tx_vec(10) => 
                           vc_write_tx_vec_10_port, vc_write_tx_vec(9) => 
                           vc_write_tx_vec_9_port, vc_write_tx_vec(8) => 
                           vc_write_tx_vec_8_port, vc_write_tx_vec(7) => 
                           vc_write_tx_vec_7_port, vc_write_tx_vec(6) => 
                           vc_write_tx_vec_6_port, vc_write_tx_vec(5) => 
                           vc_write_tx_vec_5_port, vc_write_tx_vec(4) => 
                           vc_write_tx_vec_4_port, vc_write_tx_vec(3) => 
                           vc_write_tx_vec_3_port, vc_write_tx_vec(2) => 
                           vc_write_tx_vec_2_port, vc_write_tx_vec(1) => 
                           vc_write_tx_vec_1_port, vc_write_tx_vec(0) => 
                           vc_write_tx_vec_0_port);

end SYN_structural;
